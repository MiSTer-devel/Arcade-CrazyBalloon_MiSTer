library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity SAMPLE is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(15 downto 0);
	data : out std_logic_vector(15 downto 0)
);
end entity;

architecture prom of SAMPLE is
	type rom is array(0 to  35134) of std_logic_vector(15 downto 0);
	signal rom_data: rom := (
		X"FF50",X"FEE7",X"FF03",X"FF10",X"FF33",X"FEEB",X"FEDA",X"FF07",X"FEFB",X"FF07",X"FEFD",X"FEEE",X"FF05",X"FF40",X"FF6B",X"FF82",
		X"FF7D",X"FF8E",X"FFBB",X"FFC8",X"FF7D",X"FF85",X"FF27",X"FF52",X"FF0E",X"FF78",X"FF2C",X"FF81",X"FF64",X"FF9C",X"FFC2",X"FFE5",
		X"004C",X"FFB4",X"008E",X"FFD0",X"0089",X"FF36",X"0083",X"FF1A",X"000F",X"FEF1",X"FFEF",X"FF36",X"0008",X"0013",X"0054",X"00C7",
		X"004C",X"0117",X"0079",X"00ED",X"0065",X"00C8",X"0050",X"0049",X"FF9C",X"00A6",X"FF3C",X"00CE",X"FE9D",X"013E",X"FED8",X"00EA",
		X"FFA2",X"013D",X"003A",X"00C7",X"009A",X"007C",X"01B7",X"FFD6",X"022B",X"FF36",X"0190",X"FF62",X"00CB",X"000B",X"0014",X"FFEE",
		X"002D",X"FFA4",X"00E0",X"FFE3",X"007D",X"00B9",X"FFE6",X"0195",X"FFF6",X"0107",X"00DC",X"FFDB",X"014C",X"0042",X"FFC1",X"0199",
		X"FF34",X"0125",X"FFFB",X"FFB5",X"00F0",X"FF7E",X"001A",X"0060",X"FF27",X"0068",X"FFB2",X"FED6",X"01F2",X"FE50",X"002C",X"017B",
		X"FE5A",X"0195",X"00C6",X"FF78",X"0167",X"009A",X"FFF4",X"00E7",X"008D",X"FF2F",X"FFB1",X"003C",X"FE4F",X"FED2",X"FFDF",X"FDC9",
		X"FF2A",X"FF22",X"FF14",X"FFFD",X"FEB6",X"00A1",X"0080",X"FF05",X"00FC",X"0115",X"FE8D",X"000D",X"00F0",X"FF11",X"FEDA",X"0016",
		X"FFB3",X"FD6A",X"0007",X"00AE",X"FDB9",X"FF0E",X"0131",X"FE55",X"FE88",X"0190",X"FFC2",X"FE6B",X"0086",X"018F",X"FEA8",X"005B",
		X"02AF",X"FEA4",X"0030",X"02AE",X"FFB4",X"0032",X"017C",X"011B",X"FFBB",X"007E",X"01B1",X"0022",X"FF20",X"01A1",X"0173",X"FF0D",
		X"005B",X"01DB",X"00CF",X"FF1B",X"010C",X"0235",X"003E",X"FEF9",X"0245",X"01E1",X"FEA4",X"0023",X"0279",X"0139",X"FD71",X"013D",
		X"035B",X"FF0D",X"FE92",X"0383",X"0230",X"FD64",X"00C8",X"03D5",X"FEBE",X"FD58",X"030C",X"0175",X"FC65",X"FF67",X"0385",X"FE2D",
		X"FC0F",X"0216",X"0147",X"FB42",X"FE23",X"02C9",X"FE88",X"FAD5",X"0060",X"029D",X"FC9C",X"FCA6",X"0395",X"007C",X"FBDB",X"0035",
		X"0355",X"FE01",X"FC94",X"01E0",X"00E0",X"FC11",X"FDF1",X"0337",X"FEDD",X"FBC1",X"002F",X"038B",X"FE05",X"FC3C",X"01AF",X"02D6",
		X"FC94",X"FD12",X"02CE",X"015E",X"FC78",X"FDC1",X"022E",X"FF6E",X"FBCF",X"FE80",X"009F",X"FC3C",X"FB04",X"FE98",X"FF9F",X"FC18",
		X"FBED",X"FF60",X"0084",X"FE8E",X"0008",X"0134",X"0126",X"0132",X"0246",X"0148",X"00F8",X"02C2",X"02AA",X"0170",X"0175",X"033D",
		X"0301",X"02F1",X"023D",X"032F",X"0310",X"0427",X"0360",X"01BA",X"0374",X"04A2",X"0384",X"00A6",X"01E8",X"04AE",X"0394",X"FFD0",
		X"01E4",X"0518",X"0385",X"0043",X"01E3",X"04B0",X"026D",X"00A1",X"01A2",X"0292",X"0115",X"00E7",X"0133",X"005A",X"FFB6",X"0062",
		X"FF40",X"FE66",X"FF29",X"FF44",X"FDC3",X"FCE7",X"FDC9",X"FE25",X"FCC0",X"FC4A",X"FC90",X"FC26",X"FC2E",X"FB9A",X"FBBC",X"FC46",
		X"FBFB",X"FAED",X"FBB0",X"FC83",X"FBF0",X"FB93",X"FB73",X"FC48",X"FD4E",X"FBF3",X"FAE9",X"FC6B",X"FDEA",X"FCDE",X"FADB",X"FC83",
		X"FE9D",X"FD04",X"FBA7",X"FDF7",X"FF0D",X"FD7E",X"FD55",X"FE8E",X"FE85",X"FEA0",X"FF47",X"FEDC",X"FE2A",X"FE91",X"FFDB",X"FF64",
		X"FEB2",X"FF48",X"003A",X"FFDD",X"FF5B",X"FFF2",X"00EA",X"00D7",X"FF68",X"FFD8",X"01AF",X"00BA",X"0026",X"00EA",X"0169",X"00A3",
		X"004C",X"0185",X"0179",X"FFBC",X"0025",X"0221",X"0128",X"00F2",X"018A",X"02D7",X"028C",X"021B",X"0267",X"0321",X"0374",X"02CA",
		X"01BD",X"026A",X"03A6",X"0293",X"01F6",X"0282",X"038D",X"0324",X"0254",X"02C7",X"0443",X"0320",X"0277",X"034A",X"040D",X"0398",
		X"0347",X"048D",X"0427",X"0435",X"04B9",X"057B",X"04BE",X"0488",X"05CB",X"0589",X"03D1",X"03C6",X"04CF",X"04AD",X"0284",X"02F3",
		X"0473",X"0321",X"0232",X"02CD",X"039D",X"02C2",X"019E",X"021A",X"0206",X"0176",X"01C1",X"017A",X"00B5",X"00B8",X"0172",X"00BF",
		X"FFB1",X"FFE8",X"0101",X"FFE4",X"FE77",X"FEC5",X"FFD6",X"FF57",X"FDD7",X"FEA7",X"FF10",X"FE7D",X"FDA9",X"FE00",X"FE42",X"FD8D",
		X"FD0F",X"FCE4",X"FC37",X"FC4B",X"FD1E",X"FC0B",X"FB81",X"FBF1",X"FC18",X"FB45",X"FB4B",X"FAE5",X"FB10",X"FAC3",X"FAA8",X"FA59",
		X"FA64",X"FA6D",X"FA6C",X"FAE4",X"FAA1",X"FAFC",X"FB0B",X"FA9C",X"F9F9",X"FA96",X"FB0E",X"FA5C",X"F97B",X"FA4C",X"FB3B",X"FA46",
		X"FA72",X"FB75",X"FB4E",X"FB43",X"FB32",X"FC2A",X"FC4C",X"FC2D",X"FC92",X"FD08",X"FCE5",X"FDD3",X"FE8D",X"FE6A",X"FEDC",X"FF38",
		X"009B",X"FFC2",X"0012",X"0119",X"011E",X"00EF",X"0152",X"01C6",X"01D2",X"024E",X"02D1",X"02CA",X"02E5",X"0398",X"03D5",X"03BD",
		X"03BE",X"041A",X"0439",X"040B",X"0428",X"0449",X"040B",X"04BB",X"04B7",X"0526",X"04D5",X"0549",X"0545",X"0559",X"04B8",X"04E0",
		X"0587",X"04D8",X"054B",X"0613",X"0669",X"0665",X"0697",X"07DC",X"0881",X"0786",X"06B9",X"0657",X"06C2",X"0541",X"04AB",X"03CB",
		X"02BC",X"016D",X"0114",X"01D4",X"0112",X"0010",X"FFFA",X"FF9A",X"FECC",X"FF83",X"FF62",X"FDD1",X"FCDE",X"FD43",X"FD15",X"FCAB",
		X"FC3F",X"FC87",X"FC89",X"FBC5",X"FC27",X"FBD7",X"FC55",X"FCD1",X"FC40",X"FB43",X"FBD9",X"FC13",X"FB82",X"FAFB",X"FB8D",X"FB4F",
		X"FB3D",X"FA84",X"FB90",X"FBC1",X"FAF0",X"FB27",X"FB76",X"FBA4",X"FB9E",X"FB8D",X"FC31",X"FD14",X"FC52",X"FCC0",X"FD4A",X"FDD9",
		X"FDC5",X"FE9E",X"FE76",X"FF75",X"FF68",X"FFB0",X"001E",X"0078",X"00E9",X"002C",X"009D",X"00F7",X"0128",X"0194",X"0165",X"010F",
		X"0149",X"01B3",X"011F",X"01D5",X"0117",X"011D",X"014F",X"0158",X"00A1",X"005D",X"0114",X"00FC",X"0096",X"00B0",X"00BF",X"00A4",
		X"00E1",X"008E",X"0085",X"FFF5",X"FFFB",X"007E",X"FF74",X"FF72",X"FEFC",X"0004",X"FF3F",X"FFE7",X"FF9C",X"00C6",X"FFF5",X"009D",
		X"00F0",X"010A",X"0186",X"010F",X"01EA",X"0128",X"0225",X"0127",X"02AE",X"0159",X"0390",X"01BE",X"03EC",X"02AC",X"03B4",X"034A",
		X"03F5",X"0382",X"0370",X"02FB",X"03FD",X"0207",X"034F",X"02C6",X"02DD",X"0317",X"01DB",X"0365",X"0144",X"03E8",X"01B5",X"03A5",
		X"00E3",X"0447",X"00F9",X"02B8",X"0197",X"025D",X"0299",X"008D",X"026C",X"00C2",X"01EF",X"00B4",X"0052",X"FFFD",X"0027",X"FF6F",
		X"00E7",X"FE5C",X"FFC0",X"FE8F",X"FE34",X"FF38",X"FD38",X"FEAA",X"FDE0",X"FC5E",X"FEE0",X"FD06",X"FCDA",X"FE98",X"FBEE",X"FE2B",
		X"FC72",X"FD21",X"FE0F",X"FC79",X"FD92",X"FE76",X"FC00",X"FE8A",X"FD52",X"FC46",X"0037",X"FAE3",X"FE32",X"FF85",X"FB28",X"FE60",
		X"FE68",X"FCAA",X"FDC2",X"FDB5",X"FC9C",X"FCBD",X"FE2E",X"FC45",X"FBF9",X"FDB5",X"FBF7",X"FCBB",X"FD48",X"FC55",X"FD82",X"FC24",
		X"FD43",X"FE51",X"FC61",X"FEAF",X"FF1A",X"FDB5",X"FEE2",X"0090",X"FF18",X"0051",X"01A7",X"00FB",X"FFD7",X"022B",X"034D",X"FFFF",
		X"01B9",X"0440",X"010D",X"0089",X"0471",X"024E",X"013E",X"0400",X"0453",X"011A",X"031D",X"0631",X"01A8",X"01D8",X"0692",X"01F3",
		X"0236",X"04D8",X"0377",X"0260",X"03AC",X"0462",X"02DB",X"0233",X"03EB",X"0383",X"00DB",X"02E7",X"033F",X"014F",X"0089",X"0212",
		X"028B",X"0009",X"FF67",X"01B6",X"01BC",X"FE0F",X"0001",X"018F",X"0024",X"FE02",X"0035",X"027D",X"FE01",X"FDC6",X"01C5",X"0076",
		X"FAE1",X"FE1C",X"01A4",X"FC33",X"F9DF",X"00A6",X"FEE6",X"FA38",X"FD3C",X"010D",X"FC34",X"FA0D",X"00F9",X"FF8C",X"F9A2",X"FD23",
		X"016D",X"FCCC",X"F955",X"FFA3",X"0133",X"FB16",X"FB96",X"022D",X"FF6D",X"FA3C",X"FF53",X"0250",X"FC7F",X"FB5C",X"01BD",X"005F",
		X"FB67",X"FE35",X"035B",X"FE96",X"FB38",X"006E",X"02C4",X"FCCE",X"FC34",X"022D",X"0233",X"FC26",X"FCCC",X"02C3",X"00B7",X"FBB8",
		X"FE8D",X"01EA",X"FFD9",X"FC67",X"FF7F",X"0160",X"FD2E",X"FCBB",X"0051",X"FF1C",X"FBC2",X"FD2F",X"0069",X"0131",X"FDB8",X"FFEF",
		X"01A5",X"021E",X"0321",X"047D",X"02E7",X"02EF",X"051E",X"0485",X"029C",X"03A0",X"05C0",X"039E",X"0324",X"038A",X"057A",X"057E",
		X"069F",X"06AB",X"04DC",X"0603",X"08F4",X"06C5",X"04B0",X"0721",X"08A9",X"0612",X"0269",X"0607",X"092B",X"0627",X"02FC",X"05B3",
		X"07E4",X"05B1",X"0387",X"05D0",X"05CE",X"043F",X"03CD",X"0457",X"02EB",X"027F",X"03A0",X"0272",X"FFFE",X"00A8",X"01AB",X"FEA3",
		X"FD7D",X"FEAA",X"FEF2",X"FAFE",X"FAD2",X"FCD1",X"FBBE",X"FA3F",X"F9EE",X"FA2A",X"F9CD",X"F882",X"F875",X"F88F",X"F7CF",X"F6DB",
		X"F6F0",X"F5EF",X"F62A",X"F772",X"F6BF",X"F576",X"F7E3",X"F901",X"F74E",X"F5CB",X"F85C",X"FB0F",X"F7AD",X"F625",X"F8C0",X"F9C5",
		X"F7F2",X"F7AF",X"F96C",X"F9B7",X"F9B6",X"FA62",X"F9D6",X"FA71",X"FB52",X"FC70",X"FC31",X"FB5D",X"FC82",X"FD13",X"FCA6",X"FCC3",
		X"FD69",X"FE0A",X"FDA7",X"FD32",X"FE43",X"FFE5",X"FEDB",X"FE5A",X"001C",X"0078",X"FFB2",X"FF5D",X"00F8",X"00B3",X"FEFD",X"FF75",
		X"008C",X"FFB3",X"FFB4",X"0088",X"0122",X"0173",X"01C0",X"02A9",X"03BA",X"04B2",X"044D",X"043B",X"04B4",X"06A2",X"064F",X"0518",
		X"064F",X"0806",X"0682",X"063F",X"072D",X"080E",X"070D",X"066A",X"0824",X"077D",X"06AC",X"0773",X"0942",X"0887",X"081F",X"095F",
		X"0953",X"08B9",X"08DA",X"0A0A",X"09A0",X"0858",X"089D",X"094E",X"08FE",X"0766",X"07E8",X"08FC",X"06F4",X"0671",X"07E5",X"07FC",
		X"06CA",X"057E",X"0722",X"0670",X"04C4",X"04D7",X"0468",X"033D",X"0212",X"0273",X"01C9",X"0090",X"00B0",X"0176",X"00D8",X"FF64",
		X"0061",X"0191",X"0065",X"FECB",X"FF9B",X"00DF",X"FE93",X"FDDF",X"FE85",X"FE46",X"FD79",X"FCFE",X"FCEA",X"FC3C",X"FBFA",X"FBE0",
		X"FB54",X"FA36",X"FAA2",X"FA45",X"F993",X"F953",X"F905",X"F896",X"F8A6",X"F879",X"F85A",X"F811",X"F848",X"F878",X"F7D6",X"F75F",
		X"F863",X"F910",X"F79A",X"F6D7",X"F7F7",X"F85C",X"F6E3",X"F6C8",X"F7DD",X"F7EC",X"F644",X"F708",X"F836",X"F80B",X"F82B",X"F850",
		X"F932",X"F93F",X"FA12",X"FA77",X"FA79",X"FAE6",X"FB9B",X"FCEE",X"FB4C",X"FB70",X"FCCF",X"FD6E",X"FBAE",X"FC3A",X"FE08",X"FD86",
		X"FCC0",X"FDB3",X"FF0B",X"FE57",X"FF52",X"FF9E",X"0063",X"00D2",X"0152",X"01B7",X"0108",X"00D5",X"0182",X"016F",X"0092",X"0064",
		X"012D",X"0093",X"009D",X"0197",X"0223",X"01F5",X"0296",X"0339",X"03E0",X"041D",X"0416",X"052F",X"04F1",X"0463",X"051B",X"0604",
		X"05E6",X"0644",X"07A3",X"0828",X"0805",X"08A5",X"0956",X"0906",X"078A",X"07D5",X"07CB",X"0689",X"0530",X"04A0",X"045B",X"041E",
		X"044A",X"0473",X"0436",X"03DE",X"044B",X"049E",X"043D",X"04C2",X"045A",X"0349",X"0295",X"0218",X"0226",X"01D1",X"0153",X"0097",
		X"0035",X"00D3",X"0140",X"0092",X"0028",X"0073",X"0115",X"FFB9",X"FFA2",X"0077",X"0055",X"FFE3",X"FF9B",X"FFE1",X"FFD6",X"FFD9",
		X"0006",X"FF94",X"FEC3",X"FF15",X"FEC8",X"FE08",X"FEC3",X"FEB0",X"FE6D",X"FE3F",X"FEFE",X"FF12",X"FF16",X"FFB9",X"006E",X"00E5",
		X"00BF",X"013B",X"01BA",X"019F",X"01AE",X"0221",X"022E",X"0175",X"0116",X"0193",X"01B8",X"007B",X"00AC",X"0159",X"00D4",X"000C",
		X"FF32",X"FFAF",X"FF08",X"FDCE",X"FD87",X"FDB7",X"FCBF",X"FC7C",X"FC85",X"FD2F",X"FD25",X"FC30",X"FC79",X"FCA5",X"FC8D",X"FBE4",
		X"FC1F",X"FBBA",X"FAFA",X"FB03",X"FB81",X"FA42",X"FAD5",X"FA12",X"FA7D",X"F98B",X"FA87",X"FA3C",X"F9D6",X"FAEF",X"FAC2",X"FAF4",
		X"FA21",X"FCB6",X"FB16",X"FCF6",X"FBDE",X"FE5B",X"FC36",X"FE26",X"FE28",X"FF84",X"FEC0",X"FFAE",X"FFF8",X"FF61",X"FF7E",X"009F",
		X"FFCF",X"0057",X"FFD8",X"0052",X"0077",X"FF80",X"022C",X"FFA4",X"027E",X"FF23",X"0280",X"0042",X"036F",X"00D8",X"0325",X"01D5",
		X"02FD",X"03BA",X"024A",X"056E",X"028F",X"0487",X"0296",X"0363",X"0326",X"027D",X"02BE",X"02FB",X"0150",X"02FF",X"0123",X"0161",
		X"0225",X"0080",X"031C",X"0120",X"0147",X"02DC",X"0078",X"02F9",X"0295",X"00B1",X"02F8",X"00AB",X"0257",X"025F",X"0114",X"02E2",
		X"021E",X"01A7",X"0329",X"0144",X"0312",X"03C9",X"FEA7",X"0446",X"019F",X"FFE4",X"0324",X"FF2A",X"0051",X"012D",X"FF46",X"FF47",
		X"00B9",X"002C",X"FF3A",X"00C9",X"0016",X"FE91",X"0130",X"FFC0",X"FE8F",X"013F",X"FF41",X"0045",X"004F",X"FF5E",X"01E9",X"000D",
		X"FF4D",X"01FE",X"0078",X"FF7C",X"0104",X"00A9",X"FF40",X"0005",X"01EA",X"FF82",X"FF8A",X"024B",X"0027",X"FE8F",X"0226",X"01CF",
		X"FD75",X"00F3",X"0271",X"FEF0",X"FECB",X"020B",X"0096",X"FD3C",X"01A8",X"0175",X"FCA5",X"0189",X"01A4",X"FE1F",X"0049",X"00BD",
		X"FFD3",X"FEC1",X"0028",X"006B",X"FDB0",X"FE35",X"00E7",X"FE42",X"FD0B",X"FF76",X"FFAD",X"FD77",X"FD46",X"FF75",X"FEE9",X"FC21",
		X"FD1B",X"FFD7",X"FC81",X"FB10",X"FE2B",X"FF62",X"FC4C",X"FABF",X"0042",X"FEB1",X"FA8F",X"FD20",X"016F",X"FCFA",X"FAD4",X"008C",
		X"00B5",X"FAB6",X"FDC8",X"0200",X"FCF0",X"FAE9",X"00C2",X"0117",X"F9F9",X"FD0E",X"02D8",X"FD54",X"FA50",X"00A1",X"01F2",X"FC5D",
		X"FBD0",X"028A",X"FFF6",X"F9E5",X"FF18",X"0317",X"FC42",X"FBD2",X"01A3",X"0142",X"FB54",X"FE7A",X"02D2",X"FFE3",X"FC2F",X"021C",
		X"0349",X"FCF2",X"FDCB",X"0308",X"02C4",X"FBF3",X"FF00",X"045A",X"01F0",X"FC38",X"00D8",X"056E",X"00EF",X"FD57",X"0121",X"02E9",
		X"FEF5",X"FCFC",X"00F0",X"FF9A",X"FB54",X"FE24",X"0146",X"FFC2",X"FDB7",X"FF30",X"01EA",X"02A4",X"016F",X"0290",X"0296",X"0330",
		X"040B",X"04CA",X"026A",X"03EE",X"04B4",X"040C",X"0321",X"044F",X"0603",X"0589",X"0544",X"0554",X"070B",X"06D3",X"0843",X"05E4",
		X"05F3",X"07F6",X"0869",X"0582",X"0428",X"0713",X"089C",X"0606",X"03B5",X"0734",X"08EA",X"0635",X"0514",X"07A8",X"0789",X"04BB",
		X"0442",X"053F",X"043A",X"035B",X"02E6",X"0257",X"011A",X"014B",X"0193",X"FFB2",X"FF95",X"001C",X"FF21",X"FD9F",X"FCDE",X"FDF5",
		X"FD14",X"FB67",X"FB39",X"FAF6",X"FADC",X"FA38",X"F95D",X"F976",X"F972",X"F812",X"F818",X"F89B",X"F77F",X"F6EC",X"F777",X"F75D",
		X"F764",X"F7F0",X"F6D7",X"F6EF",X"F871",X"F97D",X"F810",X"F68B",X"F954",X"FA54",X"F7CC",X"F73D",X"F9D0",X"FA17",X"F984",X"F9DE",
		X"FABC",X"FAB6",X"FBA0",X"FC49",X"FB4B",X"FB13",X"FBF6",X"FC21",X"FAFC",X"FA2C",X"FB40",X"FC10",X"FB33",X"FAED",X"FBBE",X"FD57",
		X"FCCD",X"FC10",X"FDF1",X"FEA6",X"FD6A",X"FDA0",X"FE07",X"FE79",X"FE0D",X"FE48",X"FEE7",X"FEC5",X"FE3C",X"0000",X"00C3",X"0016",
		X"00FE",X"01E7",X"030C",X"029E",X"02EE",X"03EB",X"04D4",X"047C",X"04BA",X"043D",X"055C",X"059A",X"055C",X"04BE",X"04E4",X"05E5",
		X"04BE",X"043F",X"05C1",X"0659",X"04DA",X"0549",X"0713",X"077E",X"0619",X"079D",X"08A5",X"07CA",X"0896",X"099B",X"09FA",X"08DF",
		X"09CB",X"0B1B",X"0992",X"08F1",X"0A07",X"0A22",X"08C9",X"0810",X"08A8",X"08D7",X"07C2",X"0722",X"079A",X"07BC",X"06A1",X"0601",
		X"063D",X"05B8",X"058C",X"04F5",X"0470",X"03BD",X"03EE",X"0473",X"02D5",X"021B",X"02F3",X"03DC",X"01C3",X"00B6",X"0145",X"01EA",
		X"FFAE",X"FDD3",X"FE7C",X"FE9D",X"FD50",X"FCB0",X"FC70",X"FCD3",X"FC61",X"FC4A",X"FBDD",X"FB39",X"FBA4",X"FB5B",X"FA08",X"F9AE",
		X"FA21",X"F92E",X"F866",X"F7DF",X"F7EA",X"F738",X"F742",X"F732",X"F6A2",X"F62E",X"F68B",X"F6F7",X"F5F6",X"F5AC",X"F6A9",X"F71E",
		X"F595",X"F5AB",X"F75E",X"F759",X"F658",X"F5C7",X"F7B2",X"F743",X"F63D",X"F6BA",X"F7C0",X"F7A0",X"F77F",X"F843",X"F90A",X"F9C7",
		X"FA33",X"FAE6",X"FB15",X"FB33",X"FC4C",X"FCA1",X"FC31",X"FC55",X"FE2A",X"FE69",X"FD4E",X"FE93",X"FF9D",X"FFD5",X"FF1D",X"0005",
		X"009C",X"00D8",X"0115",X"00E7",X"017A",X"01BA",X"0227",X"01EB",X"023B",X"02B9",X"0259",X"035D",X"0327",X"0358",X"03F9",X"03D2",
		X"048B",X"050C",X"053C",X"05BD",X"0638",X"06A9",X"0708",X"068B",X"07A3",X"0802",X"0807",X"087C",X"091B",X"0992",X"09EC",X"0A70",
		X"0BCE",X"0BDF",X"0A89",X"0A6E",X"0AD1",X"0A23",X"0839",X"07A3",X"0736",X"0628",X"04EC",X"0538",X"04C4",X"045C",X"049C",X"050A",
		X"04A2",X"0444",X"04F6",X"041B",X"0319",X"027A",X"0207",X"01B7",X"0017",X"0050",X"00D6",X"FFE9",X"FF63",X"FF7B",X"FEEB",X"FEF5",
		X"FF21",X"FE43",X"FD48",X"FD27",X"FCFF",X"FC3E",X"FC3F",X"FC19",X"FC30",X"FB7B",X"FB46",X"FC11",X"FB96",X"FB81",X"FBDA",X"FB54",
		X"FB93",X"FBC8",X"FBDF",X"FC4D",X"FC42",X"FC17",X"FC42",X"FCB6",X"FCBB",X"FD58",X"FDFB",X"FDBD",X"FE18",X"FE55",X"FE9C",X"FE81",
		X"FEF7",X"FFA1",X"FFB1",X"FEEB",X"FF9E",X"FFBF",X"FF42",X"FF82",X"FF97",X"FF74",X"FEC2",X"FEAC",X"FEA8",X"FD87",X"FD3B",X"FDE1",
		X"FD71",X"FD45",X"FCE7",X"FD09",X"FD92",X"FD7C",X"FD6D",X"FD4C",X"FCFC",X"FD26",X"FCD2",X"FCBD",X"FC94",X"FCE4",X"FCA4",X"FBC4",
		X"FBC0",X"FCCF",X"FD0B",X"FC0D",X"FC0B",X"FCB8",X"FCFE",X"FBB6",X"FD40",X"FBDF",X"FDD4",X"FCB9",X"FE60",X"FD13",X"FE1B",X"FE22",
		X"FEE2",X"FF23",X"FF77",X"0086",X"0022",X"020F",X"019C",X"036A",X"0312",X"045C",X"0330",X"03DA",X"03E4",X"0445",X"0263",X"0405",
		X"01BA",X"0473",X"019D",X"0405",X"0305",X"0461",X"034E",X"045C",X"05C8",X"04AD",X"05C8",X"044E",X"0762",X"03B8",X"06E8",X"03CF",
		X"056D",X"0423",X"0431",X"03BE",X"0305",X"0325",X"0373",X"022F",X"02A2",X"0206",X"011D",X"0303",X"006E",X"0162",X"00A9",X"003C",
		X"0192",X"FDE8",X"004A",X"01AD",X"FE4D",X"0069",X"FE90",X"FFE0",X"00AB",X"FDDA",X"FF82",X"FF78",X"FE1F",X"FF57",X"FD30",X"FDDF",
		X"FFC5",X"FB39",X"FEEA",X"FE44",X"FAD1",X"002C",X"FC92",X"FCCE",X"FEC3",X"FCDC",X"FD09",X"FE29",X"FCF6",X"FC98",X"FE2E",X"FDAB",
		X"FBEF",X"FDA0",X"FE13",X"FBCB",X"FE22",X"FD1F",X"FDB9",X"FE09",X"FD21",X"FFD8",X"FDDB",X"FDAF",X"0081",X"FF4F",X"FDCE",X"004E",
		X"0017",X"FF5B",X"0074",X"0137",X"0016",X"0093",X"02C3",X"00E5",X"FFC2",X"0333",X"02B5",X"FF8D",X"02E4",X"036D",X"0030",X"0239",
		X"0459",X"01A2",X"0070",X"04A9",X"03D8",X"FF78",X"0476",X"04DC",X"0026",X"02EA",X"03FD",X"0291",X"0216",X"0326",X"0359",X"0126",
		X"0210",X"0342",X"00C5",X"0018",X"0305",X"0186",X"FF63",X"0063",X"025E",X"00CA",X"FE59",X"008E",X"01D9",X"FE72",X"FDCC",X"016A",
		X"000A",X"FD5B",X"FD7E",X"01F2",X"FF37",X"FB70",X"FF9A",X"0215",X"FCC2",X"FB8A",X"01A0",X"FF82",X"F9E6",X"FD94",X"01B2",X"FB00",
		X"F9EF",X"FFE2",X"FE77",X"F856",X"FC93",X"011B",X"FAA2",X"F92F",X"002D",X"FF43",X"F8F7",X"FBE3",X"0187",X"FCCD",X"F881",X"FEC1",
		X"015E",X"F9DA",X"FB46",X"017F",X"FEAD",X"F9CB",X"FEE7",X"01EF",X"FCCD",X"FB55",X"0173",X"01BD",X"FB4A",X"FDE9",X"03C9",X"0072",
		X"FB6F",X"0053",X"0463",X"FED9",X"FB80",X"0169",X"0416",X"FE92",X"FDF8",X"02BD",X"0309",X"FF10",X"FFCC",X"035C",X"00D9",X"FD58",
		X"FFEB",X"020D",X"FD91",X"FC8C",X"FF77",X"0252",X"FF6F",X"FEB7",X"01F1",X"02F0",X"02E3",X"0463",X"048D",X"0353",X"049F",X"0589",
		X"044C",X"03B7",X"05A6",X"0640",X"0583",X"0504",X"0675",X"0763",X"07CE",X"08E8",X"0707",X"0664",X"0907",X"0901",X"05D8",X"0597",
		X"086F",X"0796",X"02E5",X"0306",X"07A4",X"07D4",X"0308",X"03C3",X"0683",X"0690",X"038A",X"0448",X"05F8",X"041C",X"02ED",X"02E0",
		X"0386",X"01B4",X"028F",X"0201",X"FF88",X"FECA",X"0093",X"FF38",X"FCB9",X"FD82",X"FE6E",X"FC16",X"F96B",X"FB43",X"FAEC",X"F9A5",
		X"F8ED",X"F8D3",X"F85A",X"F767",X"F730",X"F77A",X"F73F",X"F6B2",X"F692",X"F58F",X"F575",X"F680",X"F746",X"F57A",X"F5E0",X"F7ED",
		X"F80B",X"F5FE",X"F638",X"F9C4",X"F964",X"F64A",X"F696",X"F985",X"F881",X"F728",X"F858",X"F93A",X"F92D",X"F8FD",X"FA34",X"F9FA",
		X"FAC2",X"FB83",X"FC81",X"FB03",X"FAD4",X"FC05",X"FBD3",X"FB29",X"FB50",X"FCF0",X"FC90",X"FC0C",X"FD07",X"FEFA",X"FF55",X"FE88",
		X"FF8F",X"00F3",X"00DA",X"000D",X"011B",X"0207",X"0130",X"0056",X"01F9",X"02AD",X"01AF",X"02DF",X"03B3",X"0428",X"0360",X"04AA",
		X"0587",X"05EB",X"05D3",X"056F",X"04E9",X"062F",X"0664",X"058A",X"0596",X"0744",X"077E",X"05C9",X"067E",X"083E",X"07FA",X"0662",
		X"078D",X"0818",X"0793",X"0738",X"0944",X"0931",X"07B7",X"08CF",X"0993",X"095F",X"08BB",X"0A29",X"0AAF",X"0918",X"0894",X"09AC",
		X"0961",X"0865",X"0796",X"0836",X"0867",X"06FA",X"06EE",X"07DC",X"077B",X"064B",X"0667",X"06AA",X"0614",X"04F6",X"0530",X"03DD",
		X"02DA",X"031D",X"033E",X"014C",X"00ED",X"023C",X"0218",X"0015",X"FFA5",X"0182",X"0119",X"FF19",X"FEED",X"003F",X"FF05",X"FDB0",
		X"FDA7",X"FD34",X"FCF7",X"FC68",X"FBDF",X"FB73",X"FB18",X"FB9C",X"FAA7",X"F9C3",X"FA0D",X"FA82",X"F97A",X"F8B5",X"F8EE",X"F880",
		X"F7DB",X"F7EF",X"F73B",X"F6EC",X"F6F8",X"F6DF",X"F6BC",X"F66E",X"F660",X"F722",X"F6F1",X"F5BE",X"F68F",X"F7B4",X"F73E",X"F617",
		X"F6BB",X"F837",X"F737",X"F5E6",X"F7C7",X"F7FF",X"F794",X"F7F3",X"F8D3",X"F971",X"F99F",X"F9E0",X"FA90",X"FACF",X"FB48",X"FC79",
		X"FBF3",X"FB6F",X"FC3A",X"FCBE",X"FC97",X"FBCA",X"FC54",X"FCF3",X"FC9A",X"FCEC",X"FD90",X"FDBA",X"FE63",X"FFB8",X"FFEA",X"0069",
		X"00C8",X"0112",X"0112",X"00ED",X"0176",X"01DF",X"0153",X"00B4",X"0138",X"0224",X"0272",X"0334",X"03C4",X"03E1",X"04B3",X"05A9",
		X"0606",X"0669",X"069D",X"06A7",X"06FE",X"06AD",X"0726",X"0739",X"0851",X"08B5",X"08BE",X"09EB",X"0A56",X"0A7D",X"0B13",X"0B70",
		X"0AC2",X"091E",X"0913",X"08ED",X"07C3",X"0613",X"05D6",X"05D6",X"053A",X"055A",X"04F9",X"051E",X"04CD",X"053F",X"0492",X"04C0",
		X"04EB",X"0450",X"036D",X"0213",X"024B",X"0259",X"00FF",X"0052",X"0038",X"FFA3",X"FF6A",X"FF05",X"FEF0",X"FF1C",X"FF9F",X"FED5",
		X"FDC6",X"FE03",X"FE67",X"FE62",X"FE07",X"FDBC",X"FD3C",X"FD3D",X"FD18",X"FDD2",X"FD39",X"FCB2",X"FCE5",X"FC59",X"FC59",X"FCE9",
		X"FCFA",X"FD05",X"FD43",X"FDBE",X"FD3C",X"FD41",X"FE34",X"FE7C",X"FDB4",X"FE24",X"FE9D",X"FEA9",X"FE60",X"FF6D",X"FF82",X"FF3E",
		X"FF10",X"FF0E",X"001F",X"FF72",X"FF9D",X"0006",X"FFA7",X"FF3A",X"FEBA",X"FEE3",X"FF28",X"FE11",X"FDA9",X"FD9D",X"FD1B",X"FD71",
		X"FD70",X"FCF3",X"FCF8",X"FCFB",X"FC35",X"FB88",X"FBA3",X"FB7F",X"FBEE",X"FABD",X"FA48",X"FB0D",X"FAD1",X"FB26",X"FA7B",X"FB22",
		X"FAC8",X"FB52",X"FA38",X"FB27",X"FA8E",X"FBA9",X"FB4C",X"FC0A",X"FBA9",X"FC92",X"FDA2",X"FCEC",X"FE27",X"FDED",X"FF73",X"FE12",
		X"00F8",X"FFDE",X"01C5",X"010F",X"02DD",X"01E4",X"028C",X"02A8",X"0331",X"01B9",X"037D",X"01CF",X"03A6",X"0297",X"0351",X"03FF",
		X"03D2",X"04F1",X"03F1",X"0553",X"0366",X"068E",X"0377",X"06D3",X"036C",X"06DF",X"03F6",X"05BF",X"066C",X"04FB",X"0635",X"042D",
		X"058A",X"045D",X"03DE",X"0400",X"037D",X"01BF",X"03AC",X"00F4",X"02AD",X"0149",X"017C",X"02FB",X"00B3",X"0205",X"02AB",X"0095",
		X"02F3",X"0116",X"0102",X"021D",X"FFCD",X"0211",X"0018",X"003F",X"0152",X"FFF3",X"FFEE",X"017A",X"FEA2",X"01D8",X"FFB4",X"FE91",
		X"0361",X"FDE6",X"FFD5",X"01A2",X"FDEB",X"FF9B",X"FFA0",X"FD68",X"FDCE",X"FE6A",X"FD47",X"FCD2",X"FDB4",X"FCED",X"FCD6",X"FEDE",
		X"FD38",X"FDA4",X"FF0A",X"FD3B",X"FF56",X"FD94",X"FE2C",X"FF97",X"FC72",X"FE57",X"FF99",X"FD29",X"FD83",X"FF22",X"FDBC",X"FD13",
		X"FE87",X"FFA0",X"FD63",X"FF0F",X"00EC",X"FDE9",X"FE94",X"01BB",X"FF9F",X"FD6B",X"0188",X"006A",X"FD20",X"FFCB",X"024B",X"FE81",
		X"FD7F",X"02B8",X"FF7E",X"FD0A",X"0204",X"FF98",X"FD41",X"FFB8",X"FF42",X"FE76",X"FE4A",X"FF66",X"FE93",X"FC8E",X"FF46",X"0093",
		X"FD12",X"FDC7",X"00B0",X"0062",X"FE5F",X"FFA0",X"023E",X"FFF1",X"FDD9",X"009D",X"01F4",X"FDDA",X"FE82",X"00CB",X"0115",X"FD62",
		X"FEA0",X"0358",X"0044",X"FD4F",X"01DD",X"049B",X"FF23",X"FEEB",X"048B",X"025A",X"FDBA",X"0214",X"03BC",X"FDD8",X"FDB9",X"03EC",
		X"00B8",X"FAE1",X"00DE",X"0415",X"FD61",X"FDC6",X"047F",X"037A",X"FD98",X"0139",X"0661",X"013F",X"FD87",X"045E",X"0466",X"FDBB",
		X"FF60",X"03E8",X"00D6",X"FC03",X"0128",X"02EB",X"FE72",X"FD17",X"031A",X"018F",X"FCA5",X"FECE",X"03C5",X"FFEA",X"FB48",X"FF47",
		X"02D7",X"FDDE",X"FAD0",X"016C",X"033C",X"FDB1",X"FCF4",X"0223",X"015E",X"FC99",X"FD3B",X"00EA",X"FCBD",X"F97F",X"FC97",X"FF1C",
		X"FBFA",X"FB23",X"FD03",X"FFF4",X"FECC",X"FF53",X"00E3",X"00D7",X"0185",X"02CC",X"024F",X"00CA",X"027F",X"0359",X"0216",X"009D",
		X"0326",X"037E",X"0388",X"02E3",X"039C",X"0468",X"04C7",X"0559",X"0399",X"0477",X"0690",X"066C",X"0380",X"03AA",X"06C8",X"07C8",
		X"0445",X"03AA",X"06DA",X"0775",X"0425",X"034F",X"05E0",X"0592",X"0315",X"0281",X"0407",X"03CD",X"02B8",X"027B",X"0267",X"015C",
		X"0199",X"0085",X"FF9B",X"FF9F",X"FF74",X"FED6",X"FD63",X"FCFE",X"FD85",X"FC6C",X"FBBE",X"FB60",X"FB16",X"FB1D",X"FA58",X"F9C3",
		X"F9E9",X"FA78",X"F91A",X"F904",X"F975",X"F8D7",X"F917",X"F8C8",X"F90A",X"F976",X"F944",X"F83E",X"F908",X"FA4A",X"FAC4",X"F8F2",
		X"F7F7",X"FAF5",X"FAAE",X"F875",X"F87E",X"FB3B",X"FABC",X"FA20",X"FADA",X"FBB3",X"FB6C",X"FBF9",X"FC80",X"FBF3",X"FC41",X"FD46",
		X"FDA4",X"FBE1",X"FC2E",X"FD4A",X"FD59",X"FCC4",X"FC9D",X"FD4D",X"FE16",X"FE22",X"FD40",X"FEBD",X"FF71",X"FE88",X"FEA7",X"FF20",
		X"FF03",X"FE39",X"FE8B",X"FF2B",X"FEDC",X"FDB8",X"FFF3",X"FFB4",X"FF22",X"001D",X"016B",X"01E8",X"00EE",X"00BD",X"01FF",X"02C6",
		X"02BC",X"0254",X"0267",X"03DD",X"043A",X"045B",X"03EC",X"0560",X"05EA",X"04C5",X"0549",X"06C3",X"0680",X"05B8",X"06F8",X"083B",
		X"07E7",X"0707",X"099A",X"0959",X"086C",X"095F",X"09E1",X"0979",X"0858",X"09DD",X"0A04",X"08A6",X"07FE",X"0864",X"0842",X"0789",
		X"0726",X"0894",X"0811",X"0696",X"069B",X"077E",X"0746",X"05DF",X"0602",X"05D3",X"055E",X"04E7",X"04E6",X"043F",X"0379",X"0471",
		X"046F",X"02AF",X"020A",X"0400",X"0440",X"0143",X"00E8",X"0269",X"01E1",X"FF43",X"FECD",X"0072",X"FF46",X"FDB6",X"FE1D",X"FE5D",
		X"FDBD",X"FCF4",X"FCED",X"FC84",X"FBC4",X"FC7A",X"FBB8",X"FA8D",X"F9D7",X"FA28",X"F9A5",X"F861",X"F887",X"F82D",X"F811",X"F7B9",
		X"F7D5",X"F7B9",X"F7FE",X"F7E7",X"F815",X"F74B",X"F740",X"F824",X"F7AC",X"F626",X"F6A4",X"F737",X"F6FC",X"F5AB",X"F64B",X"F832",
		X"F695",X"F62B",X"F7D7",X"F86D",X"F7BF",X"F765",X"F84F",X"F8EF",X"F8A2",X"F98C",X"FA6D",X"F9AA",X"FA47",X"FBB6",X"FB1B",X"FB2C",
		X"FBF4",X"FDE3",X"FCCA",X"FC5C",X"FD88",X"FE4E",X"FDFF",X"FDF5",X"FED6",X"FF32",X"FFCF",X"FFF4",X"00A0",X"0155",X"0191",X"019E",
		X"01D8",X"0253",X"0263",X"02A0",X"0358",X"02E5",X"02E2",X"03B8",X"03C4",X"03FC",X"03DA",X"040B",X"0481",X"0462",X"04A2",X"049B",
		X"0485",X"0548",X"0571",X"0610",X"0761",X"084A",X"0943",X"09B1",X"0A32",X"0BAF",X"0BA4",X"0A8E",X"0A73",X"0B11",X"0A49",X"08BF",
		X"083B",X"07C0",X"06F4",X"05E6",X"058C",X"04F7",X"0516",X"04E0",X"04EA",X"040A",X"04C6",X"0471",X"0386",X"0311",X"02A2",X"023F",
		X"00F3",X"0039",X"008E",X"00E4",X"FFCB",X"FFC3",X"FF6F",X"FFFD",X"0063",X"001A",X"FFEE",X"FFD8",X"FF9E",X"FF36",X"FE7C",X"FE87",
		X"FDC8",X"FDC9",X"FD0E",X"FD20",X"FDE2",X"FD37",X"FD37",X"FD3A",X"FC75",X"FCC1",X"FCE2",X"FC93",X"FD2A",X"FCB9",X"FC8E",X"FCA1",
		X"FD34",X"FCDB",X"FD5C",X"FDE8",X"FE5E",X"FE69",X"FE92",X"FF1F",X"FF70",X"FFAB",X"FF8D",X"FF89",X"0035",X"FFEC",X"0023",X"009C",
		X"017C",X"004A",X"FFE3",X"FFC7",X"FF76",X"FED9",X"FE1E",X"FE3C",X"FE29",X"FD8E",X"FD7C",X"FD57",X"FCDB",X"FD81",X"FD73",X"FD30",
		X"FC0C",X"FCBE",X"FBE9",X"FB69",X"FAD5",X"FA7B",X"FB87",X"FA67",X"FA42",X"FA3C",X"FAB6",X"FA78",X"FB73",X"FB8C",X"FC01",X"FB2D",
		X"FC6D",X"FCA6",X"FC54",X"FD9D",X"FD2E",X"FDD5",X"FC78",X"FE65",X"FD82",X"FEE8",X"FD8B",X"FF38",X"FE45",X"0006",X"FFC1",X"009C",
		X"00A3",X"01CB",X"0233",X"026B",X"0209",X"040E",X"0238",X"0307",X"02ED",X"025D",X"038D",X"01BA",X"0440",X"01F4",X"0465",X"0173",
		X"051B",X"0299",X"05C3",X"0323",X"04E3",X"0408",X"0440",X"058F",X"02AA",X"058D",X"038F",X"0488",X"032E",X"0317",X"039D",X"031C",
		X"01BD",X"0321",X"0029",X"0208",X"0198",X"00F7",X"01EF",X"FF8A",X"019C",X"01D5",X"FF24",X"0225",X"0051",X"0049",X"019A",X"FF1A",
		X"01B0",X"FF3E",X"FFBC",X"00CF",X"FF29",X"FF7A",X"001A",X"FEB2",X"00DF",X"FEC0",X"FD95",X"0203",X"FC6D",X"FED5",X"00A4",X"FBFB",
		X"001C",X"FE87",X"FCCE",X"FEFC",X"FF0A",X"FDAF",X"FEEB",X"FFE9",X"FE2E",X"FEAA",X"FF9E",X"FD51",X"FDC2",X"FF01",X"FCFA",X"FF05",
		X"FD8B",X"FE96",X"FF99",X"FD47",X"0011",X"00CF",X"FEAC",X"FFDB",X"010F",X"FF5A",X"0043",X"0121",X"004C",X"FF4D",X"0126",X"0198",
		X"FF0E",X"010F",X"02E7",X"FFA3",X"0017",X"0347",X"FFBD",X"FF66",X"02A4",X"018F",X"FED0",X"01E7",X"0452",X"FFCA",X"00EA",X"0562",
		X"0130",X"0128",X"0462",X"01CC",X"0134",X"01F7",X"0218",X"0078",X"004E",X"026C",X"0143",X"FE70",X"011E",X"0232",X"FF13",X"FEFA",
		X"0169",X"00CC",X"FE81",X"FF61",X"017A",X"006B",X"FD68",X"00D4",X"0175",X"FEF3",X"FE2B",X"00F3",X"01C8",X"FB86",X"FDD3",X"01E0",
		X"FF29",X"FA91",X"FF4E",X"0208",X"FC45",X"FBD6",X"0216",X"FF9B",X"FA71",X"FF59",X"00FF",X"FB57",X"FAC7",X"01F3",X"FEB7",X"F8F2",
		X"FEF7",X"027D",X"FC17",X"FA70",X"0199",X"011A",X"FA41",X"FCAE",X"01BE",X"FCF8",X"F8C9",X"FF4B",X"006E",X"FA0B",X"FB49",X"0180",
		X"FDDD",X"F9FF",X"FEB2",X"01F9",X"FC30",X"FA7D",X"0153",X"0069",X"FA8A",X"FBE2",X"025D",X"FF5F",X"FA5E",X"FE0E",X"0330",X"FF0D",
		X"FBB0",X"012C",X"03C7",X"FF5C",X"FD18",X"01CF",X"01B5",X"FDA9",X"FD61",X"01A8",X"FE2F",X"FB14",X"FE7E",X"0190",X"008C",X"FDFD",
		X"0011",X"02A9",X"0297",X"0359",X"044A",X"02B4",X"0370",X"04FF",X"04BC",X"0310",X"0583",X"065D",X"0565",X"04A1",X"0665",X"0863",
		X"08B8",X"0924",X"085D",X"080D",X"09AA",X"0AB5",X"082C",X"0744",X"08E5",X"09E9",X"0601",X"0543",X"087F",X"0A39",X"070D",X"0518",
		X"0872",X"0957",X"067C",X"05C7",X"07E8",X"064C",X"04C9",X"03E4",X"0495",X"03CD",X"037C",X"0458",X"0267",X"00DD",X"015E",X"0140",
		X"FFB2",X"FEFA",X"FF79",X"FE5D",X"FB6D",X"FBE1",X"FCA9",X"FB54",X"FA26",X"F94A",X"F8FC",X"F915",X"F7DC",X"F7DD",X"F847",X"F7B3",
		X"F681",X"F620",X"F679",X"F5BB",X"F6C9",X"F6EB",X"F5BA",X"F748",X"F772",X"F5F0",X"F542",X"F77D",X"F90A",X"F584",X"F494",X"F78B",
		X"F78B",X"F508",X"F5F9",X"F7D8",X"F7D3",X"F7AA",X"F89A",X"F814",X"F843",X"FA6A",X"FB0A",X"F9CD",X"F8CD",X"FA89",X"FAD5",X"FA13",
		X"F965",X"FB4B",X"FBAA",X"FAEC",X"FAF1",X"FC32",X"FD91",X"FC21",X"FC81",X"FE14",X"FD51",X"FD87",X"FE46",X"FEFA",X"FE78",X"FDC9",
		X"FE9A",X"FF6B",X"FE5B",X"FE62",X"0038",X"0024",X"008F",X"00CF",X"02D3",X"0386",X"035E",X"034B",X"0446",X"055F",X"056D",X"0513",
		X"0514",X"05DE",X"05B2",X"0519",X"053E",X"0641",X"0701",X"0627",X"066E",X"07B5",X"07A6",X"070E",X"07F7",X"092B",X"07D5",X"0799",
		X"0918",X"08C5",X"0854",X"0938",X"0A00",X"099A",X"08F2",X"0A5F",X"0B0B",X"0A3E",X"0A2D",X"0B25",X"0BD4",X"0A88",X"0A0B",X"0B0C",
		X"0B5B",X"098A",X"09AB",X"0A13",X"0977",X"087F",X"084F",X"0854",X"0748",X"075E",X"0767",X"064C",X"0538",X"061D",X"068D",X"051E",
		X"03B0",X"0481",X"056B",X"03BB",X"01F5",X"02AF",X"02E9",X"007B",X"FFED",X"FFEE",X"0004",X"FF49",X"FDEA",X"FE51",X"FD84",X"FD41",
		X"FCFE",X"FBB5",X"FAEF",X"FB7E",X"FAC1",X"F9CC",X"F99E",X"F9DF",X"F9AC",X"F964",X"F8FB",X"F8D1",X"F83C",X"F836",X"F80D",X"F742",
		X"F680",X"F679",X"F637",X"F50D",X"F4DA",X"F5F4",X"F5B3",X"F3E4",X"F385",X"F4E4",X"F5CA",X"F35F",X"F497",X"F634",X"F529",X"F4B7",
		X"F5DB",X"F6E2",X"F6AF",X"F71B",X"F7DB",X"F849",X"F7E0",X"F8F7",X"F958",X"F881",X"F964",X"F9E9",X"FA58",X"F928",X"FA0A",X"FB7E",
		X"FB56",X"FB19",X"FBD6",X"FD12",X"FD0F",X"FD93",X"FDD6",X"FEA5",X"FEBB",X"FECA",X"FF06",X"FEFE",X"FF89",X"FFCD",X"FFDE",X"0073",
		X"0070",X"0147",X"0175",X"01EE",X"0230",X"02C4",X"0392",X"03D8",X"03F8",X"0415",X"041F",X"0409",X"04DE",X"0479",X"04A0",X"0537",
		X"05DA",X"0683",X"074C",X"083A",X"0993",X"09DA",X"0AB7",X"0BDC",X"0B74",X"09C8",X"09E4",X"0A5F",X"08D7",X"0739",X"069F",X"0705",
		X"0656",X"06B7",X"06B5",X"0700",X"0661",X"0678",X"063E",X"055F",X"0580",X"04A3",X"03EF",X"027C",X"01F3",X"0238",X"0119",X"0091",
		X"013A",X"00E0",X"00B2",X"0102",X"0149",X"01A6",X"01F9",X"016B",X"006D",X"0056",X"0079",X"FFA9",X"FF69",X"FEC7",X"FED4",X"FE81",
		X"FE0B",X"FEA9",X"FEF2",X"FE2B",X"FE1D",X"FEB3",X"FE1F",X"FE61",X"FEA1",X"FF14",X"FECB",X"FE74",X"FEE2",X"FEF7",X"FEBD",X"FF5F",
		X"FFA8",X"FF95",X"FFAA",X"FFC0",X"0086",X"0058",X"0071",X"00F7",X"00B2",X"00C9",X"00AB",X"0130",X"002B",X"FFBC",X"0000",X"FF92",
		X"FE84",X"FDE1",X"FE96",X"FE36",X"FDB0",X"FD64",X"FE2A",X"FD55",X"FD26",X"FD11",X"FD1C",X"FCBC",X"FC4C",X"FC09",X"FBCF",X"FBD4",
		X"FADF",X"FBC0",X"FAD0",X"FA9E",X"FADD",X"FAC0",X"FA4F",X"FA59",X"FB11",X"FAF3",X"FAFC",X"F9E4",X"FB58",X"F9F0",X"FC16",X"FAB0",
		X"FBBF",X"FAA1",X"FC5D",X"FC75",X"FC97",X"FCA2",X"FD1A",X"FD6D",X"FD36",X"FECE",X"FDFC",X"FF93",X"FE31",X"0014",X"FEDF",X"0074",
		X"0028",X"FFE3",X"FFD1",X"01AF",X"FF20",X"01A0",X"FF4E",X"0238",X"004A",X"0187",X"00BB",X"01FB",X"019C",X"015F",X"02E8",X"0205",
		X"052C",X"0199",X"05F4",X"02CF",X"062B",X"042A",X"04B8",X"044F",X"036A",X"0435",X"03C7",X"033F",X"03F0",X"02D2",X"02FB",X"03F1",
		X"01DB",X"0414",X"018F",X"02BE",X"0288",X"00E8",X"031E",X"019B",X"00C2",X"036C",X"0027",X"0273",X"019B",X"00E1",X"0331",X"007C",
		X"01FE",X"0274",X"0197",X"024D",X"01D9",X"00AC",X"0459",X"FFF5",X"0130",X"03FB",X"FE64",X"0224",X"0195",X"FF0A",X"01DC",X"00BD",
		X"FFC0",X"00F2",X"012C",X"FF77",X"003E",X"00C3",X"FE9B",X"FF8C",X"00CB",X"FEDC",X"FFE1",X"FF9C",X"FF12",X"00CD",X"FE7A",X"00B8",
		X"002D",X"FDC1",X"0038",X"FFBF",X"FDF4",X"FF07",X"0000",X"FE98",X"FE97",X"0000",X"FFD1",X"FDA7",X"005E",X"0130",X"FDE4",X"004C",
		X"0265",X"FE99",X"FFC0",X"039D",X"0020",X"FEBB",X"022C",X"0246",X"FEB0",X"00BE",X"0417",X"FE8E",X"FFC8",X"035A",X"FF3F",X"FFD3",
		X"00E3",X"FFE3",X"FEE6",X"FEEB",X"FF79",X"FDB2",X"FCE3",X"FF5E",X"FE96",X"FBCA",X"FDAF",X"FF85",X"FD8B",X"FC3F",X"FE6D",X"FF88",
		X"FD4F",X"FC9C",X"FFE8",X"FEBA",X"FB98",X"FE2A",X"FFC2",X"FE3C",X"FB14",X"FF2B",X"010A",X"FC1D",X"FC0D",X"013E",X"00B1",X"FAED",
		X"FE82",X"0353",X"FD96",X"FBF6",X"0217",X"FFF1",X"FAC4",X"FD96",X"01D7",X"FBC4",X"F9B9",X"0148",X"FFCE",X"F983",X"FDAB",X"02C2",
		X"FE33",X"FA68",X"011C",X"02DF",X"FBCA",X"FBC5",X"0348",X"FF82",X"FA64",X"FF27",X"0265",X"FCC7",X"FC33",X"0318",X"01F9",X"FD3F",
		X"002A",X"05F3",X"00CE",X"FDD1",X"02C4",X"0595",X"FED0",X"FD64",X"0367",X"03A3",X"FD03",X"FDFC",X"0489",X"0311",X"FE31",X"0070",
		X"04DB",X"0134",X"FD80",X"00B5",X"0232",X"FC75",X"FB9B",X"0033",X"FF8A",X"FC88",X"FD86",X"00C2",X"0198",X"0046",X"020B",X"02F7",
		X"0368",X"0457",X"0546",X"0390",X"03CD",X"05C4",X"0567",X"03F3",X"041A",X"05FE",X"05DB",X"05D0",X"04CF",X"05E4",X"0666",X"0724",
		X"052D",X"048B",X"0669",X"0740",X"0536",X"02C3",X"0506",X"0716",X"05A6",X"01D2",X"03D2",X"0708",X"050E",X"0201",X"0399",X"0584",
		X"0350",X"0164",X"01EC",X"02E2",X"01F8",X"00A2",X"014B",X"0141",X"00DC",X"00FC",X"000D",X"FF20",X"FF18",X"FF07",X"FD59",X"FC37",
		X"FC4E",X"FC83",X"FA90",X"FA4A",X"FAEA",X"FA78",X"FA20",X"F903",X"F91C",X"F90A",X"F82C",X"F6AF",X"F6BB",X"F64A",X"F5C1",X"F59E",
		X"F576",X"F60B",X"F72B",X"F6B5",X"F63A",X"F805",X"F8DF",X"F856",X"F622",X"F7E8",X"FA24",X"F80B",X"F656",X"F895",X"FA78",X"F911",
		X"F93D",X"F9DF",X"FABC",X"FB95",X"FC05",X"FBEA",X"FB9D",X"FC4B",X"FDAE",X"FCCD",X"FBDD",X"FD71",X"FDF7",X"FDCD",X"FD6B",X"FE3B",
		X"FEDA",X"FF15",X"FF48",X"FFB6",X"013C",X"0056",X"0044",X"010C",X"012F",X"0113",X"0073",X"00CF",X"011F",X"0008",X"0091",X"029E",
		X"0202",X"022D",X"0348",X"050A",X"0512",X"0517",X"0575",X"0650",X"06F5",X"0653",X"05CC",X"0637",X"075F",X"06CD",X"0697",X"073A",
		X"08EA",X"0866",X"074C",X"07EC",X"092F",X"07CB",X"06A9",X"0817",X"0871",X"0703",X"0745",X"095B",X"0889",X"081C",X"096A",X"0A19",
		X"08FE",X"08AA",X"09A7",X"08A7",X"0746",X"06F2",X"0729",X"0708",X"05AE",X"05CC",X"06C9",X"05F1",X"0540",X"05D2",X"0671",X"05C7",
		X"0481",X"04C9",X"0516",X"03B1",X"0387",X"0361",X"023F",X"01AE",X"029E",X"01A7",X"FFDB",X"000B",X"00BB",X"FF82",X"FD9B",X"FE84",
		X"FEFC",X"FDAF",X"FBFA",X"FCF0",X"FD9D",X"FC8D",X"FBC8",X"FBB2",X"FBB4",X"FB5E",X"FB09",X"FADD",X"F9F7",X"FA4E",X"FACD",X"F95B",
		X"F94E",X"F954",X"F9A0",X"F88C",X"F845",X"F872",X"F800",X"F7C6",X"F7E5",X"F7B6",X"F6E4",X"F76F",X"F7C7",X"F7DB",X"F715",X"F7E6",
		X"F8D1",X"F801",X"F6D7",X"F7EC",X"F8F4",X"F76F",X"F66F",X"F7E9",X"F89D",X"F6AE",X"F724",X"F8FB",X"F8CF",X"F85E",X"F90B",X"FA3A",
		X"FA49",X"FA3E",X"FB6B",X"FB88",X"FB3B",X"FC12",X"FCFC",X"FC12",X"FC74",X"FDCD",X"FE22",X"FCCF",X"FD4B",X"FEC7",X"FEA8",X"FE55",
		X"FF3C",X"0023",X"00AD",X"010B",X"00CD",X"022B",X"027A",X"0253",X"02BF",X"0299",X"02BA",X"02DA",X"0335",X"03CA",X"033C",X"0436",
		X"0442",X"03F6",X"0498",X"04F5",X"050B",X"04FF",X"056D",X"05E7",X"0594",X"050B",X"0616",X"0695",X"069A",X"06FB",X"0847",X"08DB",
		X"08F3",X"0A53",X"0B7A",X"0B6C",X"0A5C",X"0A57",X"0A84",X"08FC",X"08BD",X"084A",X"0782",X"05EB",X"053F",X"0604",X"05BC",X"0580",
		X"0599",X"0579",X"0516",X"052F",X"04B9",X"03AC",X"0341",X"0352",X"01CB",X"0115",X"00AE",X"00B1",X"0041",X"FF23",X"FF8E",X"FEB2",
		X"FEFE",X"FF25",X"FE61",X"FE18",X"FE99",X"FEB8",X"FD58",X"FD6C",X"FDCF",X"FD94",X"FDB1",X"FDB6",X"FDF3",X"FE2E",X"FDB1",X"FE33",
		X"FDE9",X"FD70",X"FDDE",X"FD3A",X"FCCE",X"FD8F",X"FD95",X"FCF9",X"FD0E",X"FD8D",X"FCFE",X"FCCE",X"FCED",X"FDBE",X"FDD2",X"FD8B",
		X"FE63",X"FE84",X"FEEE",X"FF4D",X"FF5A",X"FFBE",X"FF2D",X"FFA0",X"FF97",X"FF50",X"FE8B",X"FEA0",X"FECC",X"FF3F",X"FE38",X"FDC4",
		X"FE6D",X"FDB1",X"FD3B",X"FD00",X"FCDB",X"FC77",X"FC92",X"FBBD",X"FBE7",X"FBC1",X"FBA0",X"FAEB",X"FAE2",X"FADD",X"FA97",X"FB0D",
		X"FAA0",X"FA30",X"FA6F",X"FB08",X"FA0F",X"FA60",X"FA03",X"FABC",X"F965",X"FB72",X"FA96",X"FB1D",X"FAC2",X"FC70",X"FB35",X"FB74",
		X"FCF2",X"FD79",X"FDBD",X"FDB2",X"0050",X"FEE0",X"0128",X"0068",X"0282",X"019E",X"0335",X"0254",X"0264",X"02A5",X"03C2",X"020F",
		X"0377",X"0248",X"04EC",X"0294",X"04B6",X"0432",X"04A1",X"044A",X"038F",X"0566",X"037D",X"058F",X"02A0",X"0689",X"0304",X"0695",
		X"03BE",X"05C1",X"054F",X"04B7",X"060D",X"0429",X"05B3",X"048F",X"043F",X"04BC",X"045B",X"02BA",X"03F7",X"01A2",X"0342",X"01DC",
		X"01EC",X"0395",X"0108",X"02BA",X"0381",X"011F",X"040F",X"0230",X"025A",X"02C5",X"0051",X"0238",X"0096",X"002E",X"00C0",X"FF71",
		X"0015",X"010C",X"FDB4",X"01AF",X"FFE2",X"FE11",X"02BE",X"FDED",X"FF73",X"00A2",X"FD9D",X"FF52",X"FF40",X"FD68",X"FDDE",X"FF6B",
		X"FDB6",X"FDA2",X"FF7E",X"FE39",X"FCDF",X"FF8A",X"FD67",X"FE0B",X"FEB6",X"FD47",X"FEF2",X"FC97",X"FD5B",X"FF28",X"FC6D",X"FCBF",
		X"FEEB",X"FCD1",X"FD8C",X"FEF9",X"FE45",X"FD33",X"FEFE",X"008B",X"FD43",X"FED4",X"0174",X"FDB3",X"FD72",X"010D",X"FF6C",X"FC31",
		X"00B1",X"0167",X"FE2C",X"FF67",X"0325",X"00E0",X"FE7C",X"0383",X"01DC",X"FEFC",X"02C2",X"00FE",X"FF35",X"00DC",X"003A",X"FEDE",
		X"FE60",X"FFBA",X"FF6E",X"FD04",X"FE5F",X"00F4",X"FE97",X"FE1F",X"FFFF",X"0044",X"FEA2",X"FF0B",X"0070",X"FFDD",X"FD6D",X"FF58",
		X"01B6",X"FEA9",X"FE8E",X"00B6",X"027E",X"FD9B",X"FDD0",X"0387",X"011F",X"FCD9",X"FFD0",X"038C",X"FDD6",X"FCB9",X"0183",X"004A",
		X"FB22",X"FF6D",X"0274",X"FCF9",X"FBEA",X"02B3",X"0158",X"FA66",X"FF7C",X"04E6",X"FE59",X"FBA9",X"0281",X"0379",X"FC49",X"FD68",
		X"03C9",X"FFF9",X"FA45",X"0052",X"03B1",X"FD6F",X"FCBF",X"02E2",X"01CD",X"FC2D",X"006B",X"03BA",X"FFD8",X"FC2F",X"022B",X"0229",
		X"FC5B",X"FC9E",X"031F",X"0121",X"FB42",X"FE66",X"041D",X"016D",X"FC22",X"01F9",X"05B9",X"016C",X"FD47",X"01F4",X"02F5",X"FDD7",
		X"FC9D",X"00B2",X"FE44",X"F97F",X"FD17",X"0197",X"FFAC",X"FCA4",X"FF2F",X"02F9",X"0160",X"0157",X"03C1",X"02E9",X"0218",X"033A",
		X"03E8",X"01AF",X"02D8",X"0419",X"0333",X"01AF",X"03A1",X"05B2",X"0630",X"0476",X"04CE",X"05FB",X"0565",X"0722",X"04CA",X"0414",
		X"061D",X"06AA",X"0384",X"020D",X"054B",X"06E2",X"04B1",X"0282",X"0631",X"0713",X"04C5",X"03E9",X"05A1",X"05BE",X"032C",X"02D5",
		X"034A",X"0317",X"024E",X"02CE",X"01FD",X"008C",X"00B1",X"00AC",X"FF9C",X"FF50",X"FF9A",X"FEDE",X"FC56",X"FB26",X"FCED",X"FC05",
		X"FA86",X"FA0C",X"FA35",X"F9FA",X"F8C9",X"F8CB",X"F97F",X"F95D",X"F799",X"F82A",X"F8E4",X"F831",X"F7D1",X"F92A",X"F881",X"F9E2",
		X"F996",X"F862",X"F91C",X"F9FB",X"FB77",X"F875",X"F7CE",X"F9A3",X"FA66",X"F83F",X"F8F2",X"FAC4",X"F9EE",X"F986",X"F9FC",X"FAA9",
		X"F9C5",X"FB62",X"FBE9",X"FAF4",X"FA93",X"FC07",X"FCD9",X"FBCD",X"FB78",X"FCAC",X"FD9C",X"FC9B",X"FCB4",X"FDF1",X"FEEC",X"FE2C",
		X"FD30",X"FF6A",X"FF46",X"FE7B",X"FF39",X"002C",X"FFB8",X"FF64",X"0033",X"010F",X"00C2",X"FF63",X"0233",X"024F",X"0125",X"01D5",
		X"03C8",X"03F0",X"02A1",X"02AC",X"03D6",X"0453",X"0424",X"03CB",X"0426",X"0566",X"056D",X"0488",X"04D2",X"05F1",X"066D",X"04E3",
		X"04FD",X"06B2",X"0754",X"05E2",X"0626",X"07E9",X"07DD",X"0661",X"07F6",X"0890",X"0785",X"07E0",X"08ED",X"0908",X"0746",X"08CE",
		X"0972",X"084D",X"0774",X"085E",X"0899",X"0684",X"063A",X"0788",X"07F3",X"065F",X"05EC",X"0747",X"070E",X"05C0",X"05BA",X"0605",
		X"04F5",X"04CA",X"0447",X"040C",X"026D",X"0351",X"03CD",X"028C",X"015E",X"022E",X"037C",X"01A5",X"FFFA",X"00BD",X"013C",X"FF1D",
		X"FDDB",X"FECB",X"FED6",X"FD81",X"FC82",X"FD05",X"FCC9",X"FC55",X"FC96",X"FBB0",X"FB50",X"FB65",X"FB32",X"FA39",X"F9DF",X"F9DB",
		X"F958",X"F912",X"F926",X"F8AD",X"F850",X"F7E4",X"F7A9",X"F72F",X"F64D",X"F62F",X"F600",X"F567",X"F49B",X"F551",X"F563",X"F3DF",
		X"F3EE",X"F560",X"F69D",X"F556",X"F557",X"F7B7",X"F74F",X"F667",X"F72B",X"F836",X"F835",X"F83B",X"F93B",X"F9E9",X"F9F5",X"FA79",
		X"FB91",X"FB21",X"FBE9",X"FCCD",X"FCBC",X"FC35",X"FCC2",X"FE1E",X"FE2F",X"FDE8",X"FEB8",X"FF3B",X"FF6E",X"003F",X"00B3",X"00BB",
		X"00D6",X"010D",X"00AC",X"00B1",X"019B",X"01F4",X"024E",X"02F4",X"0304",X"0368",X"03F8",X"0442",X"04E7",X"04B1",X"0499",X"04FC",
		X"0540",X"05C7",X"05F3",X"06B0",X"0733",X"06DC",X"06D1",X"080C",X"0879",X"092A",X"0974",X"09D2",X"0A68",X"0AD3",X"0B30",X"0C3F",
		X"0BC6",X"0A67",X"09B4",X"0A44",X"09D6",X"07F4",X"07A2",X"0707",X"0683",X"05C4",X"05BA",X"0594",X"0502",X"054C",X"058C",X"0412",
		X"03DA",X"0466",X"0329",X"01B4",X"00C0",X"0055",X"FF92",X"FDD2",X"FE67",X"FED3",X"FE81",X"FE6F",X"FE86",X"FF88",X"004D",X"0043",
		X"FFF8",X"FFBF",X"FF93",X"FE68",X"FD8E",X"FD73",X"FCDB",X"FC99",X"FC4F",X"FC75",X"FD1F",X"FCF5",X"FCB1",X"FCCA",X"FC6E",X"FC3D",
		X"FBA9",X"FBBE",X"FC5F",X"FC06",X"FB25",X"FB74",X"FC02",X"FB89",X"FC45",X"FCD4",X"FD39",X"FDDB",X"FEC3",X"FF15",X"FF72",X"003D",
		X"009B",X"0072",X"0069",X"008B",X"0083",X"FFE3",X"FFE7",X"FF52",X"FF21",X"FE6B",X"FE07",X"FDF8",X"FD42",X"FDB0",X"FDBD",X"FD1E",
		X"FC99",X"FCCD",X"FC3B",X"FC79",X"FBF2",X"FB64",X"FA95",X"FAA4",X"FAB4",X"FA24",X"FA14",X"F9DE",X"FAAA",X"FA92",X"F9B2",X"F9CA",
		X"FBA7",X"FAB1",X"FAC5",X"F9E7",X"FB6E",X"FAB4",X"FB18",X"FBBF",X"FB42",X"FC81",X"FCAB",X"FDB0",X"FCB4",X"FECC",X"FDB6",X"FFB7",
		X"FE4F",X"0076",X"FF3B",X"00E6",X"0023",X"005B",X"007E",X"01E3",X"01CE",X"0102",X"0167",X"0302",X"01BF",X"0202",X"024B",X"02A2",
		X"03A6",X"0254",X"04D4",X"02D6",X"0674",X"0380",X"068E",X"0397",X"071F",X"050B",X"0699",X"05FB",X"05C0",X"0759",X"04AD",X"076B",
		X"0483",X"0669",X"04CF",X"0493",X"04E7",X"04A7",X"0319",X"04D2",X"0258",X"0397",X"037B",X"02A4",X"0420",X"01A4",X"042B",X"042B",
		X"01CD",X"0428",X"02D3",X"01B7",X"02D1",X"FF91",X"027B",X"00A8",X"FFC4",X"0164",X"0058",X"011F",X"0205",X"003C",X"0356",X"01B2",
		X"FF07",X"0480",X"FF07",X"007B",X"0273",X"FDFE",X"000D",X"FF84",X"FE17",X"FF7C",X"FFF0",X"FE26",X"FF1A",X"0060",X"FE1E",X"FE6D",
		X"0000",X"FE0C",X"FD81",X"FE87",X"FC98",X"FE65",X"FCB1",X"FD04",X"FEFF",X"FBCA",X"FD03",X"FEE5",X"FC67",X"FCCF",X"FE82",X"FD42",
		X"FDBE",X"FE7C",X"FDED",X"FD06",X"FEEB",X"0047",X"FD07",X"FEF2",X"01CF",X"FE9E",X"FDCB",X"0227",X"0018",X"FDB1",X"015C",X"0105",
		X"FE62",X"FEF3",X"0221",X"FE51",X"FD5B",X"01F2",X"FDCD",X"FCB5",X"FF61",X"FDC5",X"FD31",X"FDC7",X"FEE7",X"FDC0",X"FCA9",X"FF3D",
		X"FFF5",X"FCBC",X"FE76",X"0040",X"FE25",X"FCB3",X"FED4",X"FFDF",X"FD71",X"FD2A",X"FFE5",X"0014",X"FC97",X"FF98",X"020F",X"FFC0",
		X"FDA9",X"0097",X"0382",X"FD8A",X"FDDD",X"0341",X"0292",X"FC33",X"FEDC",X"03CA",X"FE48",X"FBBC",X"01D2",X"00BA",X"FA9E",X"FE36",
		X"022F",X"FD9B",X"FB14",X"0267",X"01A1",X"FB2C",X"FF70",X"0562",X"0042",X"FCD1",X"0248",X"0460",X"FD9C",X"FD16",X"038C",X"011F",
		X"FB69",X"000D",X"03D6",X"FE96",X"FD85",X"0459",X"0376",X"FE67",X"00CE",X"0594",X"00EF",X"FCD9",X"0252",X"03B8",X"FDF9",X"FCE9",
		X"034C",X"0321",X"FD23",X"FE22",X"04A1",X"030F",X"FEA1",X"01CB",X"0585",X"0231",X"FEC2",X"01FF",X"0226",X"FDE2",X"FBEF",X"FF83",
		X"FDC0",X"F9BB",X"FB95",X"FFAA",X"001B",X"FE02",X"FFDB",X"0214",X"02CF",X"03F4",X"05A5",X"02E3",X"02E6",X"046B",X"043E",X"0156",
		X"034B",X"054B",X"03A0",X"02F4",X"03ED",X"0681",X"0645",X"07A4",X"0788",X"05E2",X"0739",X"094C",X"0711",X"045D",X"05B9",X"076C",
		X"043E",X"00A7",X"037F",X"0720",X"049D",X"01C8",X"0480",X"06AB",X"051C",X"0310",X"056F",X"0585",X"035A",X"0277",X"02A4",X"0176",
		X"0139",X"01FD",X"0022",X"FEB7",X"FF4E",X"0028",X"FDA6",X"FDD2",X"FF0A",X"FEF0",X"FB8D",X"FB5E",X"FCEE",X"FB00",X"F9B0",X"F92A",
		X"F88B",X"F727",X"F674",X"F630",X"F6E8",X"F688",X"F598",X"F5A0",X"F5BF",X"F5ED",X"F739",X"F74A",X"F5AD",X"F783",X"F850",X"F6F7",
		X"F586",X"F732",X"FA15",X"F75D",X"F5B0",X"F7BA",X"F959",X"F72F",X"F778",X"F8E8",X"F932",X"F962",X"F9D0",X"F952",X"F9E7",X"FB6B",
		X"FBD5",X"FB54",X"FA4B",X"FBE3",X"FC55",X"FBEE",X"FC24",X"FD2A",X"FD47",X"FDA6",X"FDF1",X"FEBF",X"0050",X"FFDE",X"FEFD",X"002D",
		X"FFC9",X"FFFB",X"FF67",X"00A1",X"0101",X"000F",X"0047",X"022C",X"01B6",X"0164",X"0331",X"034C",X"03C6",X"0310",X"04C5",X"05B6",
		X"0647",X"0571",X"05A8",X"06AA",X"07C5",X"078C",X"072E",X"0800",X"08B9",X"0812",X"074C",X"083C",X"092A",X"0820",X"0772",X"0879",
		X"08F1",X"07AA",X"085B",X"0AAC",X"09D6",X"08B0",X"098C",X"09E1",X"0904",X"08B8",X"09DA",X"098D",X"07CD",X"0827",X"0908",X"08AD",
		X"080C",X"0890",X"092D",X"0794",X"0725",X"0851",X"0871",X"0774",X"06FC",X"07A7",X"073C",X"060C",X"05BE",X"05E6",X"04D7",X"046D",
		X"047C",X"038F",X"01D5",X"0267",X"0335",X"01CD",X"FFD3",X"FFE3",X"00F3",X"FFBB",X"FDCF",X"FE41",X"FED3",X"FD11",X"FC43",X"FCC8",
		X"FCDA",X"FC9C",X"FBC2",X"FBCF",X"FAE9",X"FA26",X"FA69",X"F98E",X"F89C",X"F8EF",X"F917",X"F81D",X"F7B4",X"F81B",X"F7B4",X"F7C1",
		X"F72D",X"F6EB",X"F629",X"F569",X"F60E",X"F4FF",X"F3F9",X"F410",X"F4C1",X"F3C9",X"F30E",X"F478",X"F5A9",X"F496",X"F395",X"F576",
		X"F6BA",X"F4BE",X"F4C7",X"F6A5",X"F6A1",X"F56F",X"F5EE",X"F6D9",X"F6F7",X"F73F",X"F817",X"F927",X"F944",X"F9E0",X"FAB3",X"FA2B",
		X"FA93",X"FC2C",X"FCA4",X"FB97",X"FBFB",X"FDD0",X"FDA3",X"FD8C",X"FDEB",X"FEC8",X"FEFA",X"FF15",X"FF66",X"00A3",X"01D4",X"025E",
		X"02F7",X"0349",X"0393",X"03FE",X"0485",X"04D1",X"04C7",X"0510",X"056C",X"0575",X"05FB",X"0651",X"06C6",X"0742",X"0746",X"0779",
		X"0879",X"080B",X"0926",X"08F3",X"08AD",X"08CA",X"095B",X"09F1",X"09DA",X"0AA2",X"0B94",X"0BAF",X"0B36",X"0C3E",X"0CA6",X"0B3F",
		X"0AC9",X"0BFA",X"0A8F",X"094F",X"08B5",X"0893",X"07BE",X"06E7",X"06DF",X"0603",X"0535",X"054F",X"0521",X"03F5",X"03C0",X"03B3",
		X"0364",X"0211",X"0173",X"01FE",X"0152",X"FFFF",X"FF90",X"FF2E",X"FF4E",X"FEF7",X"FE4D",X"FE0E",X"FEB8",X"FF5E",X"FE1B",X"FD7D",
		X"FDDF",X"FDAC",X"FD44",X"FC9F",X"FBDB",X"FC54",X"FBC7",X"FBEC",X"FBD1",X"FB47",X"FB07",X"FAEA",X"FAAF",X"FB1F",X"FB4D",X"FBAA",
		X"FB93",X"FB93",X"FBF8",X"FC0E",X"FC03",X"FC30",X"FD02",X"FCCE",X"FCDD",X"FD20",X"FDD1",X"FDFC",X"FE86",X"FEB6",X"FE90",X"FE24",
		X"FEA4",X"FF48",X"FED8",X"FF1E",X"FE9C",X"FE2A",X"FE07",X"FD3C",X"FD89",X"FD9F",X"FCAB",X"FC63",X"FCA4",X"FC43",X"FC0B",X"FBC1",
		X"FC0C",X"FC33",X"FBBF",X"FB99",X"FB98",X"FBC9",X"FB84",X"FC32",X"FBD1",X"FBD8",X"FC27",X"FC4E",X"FBE6",X"FB80",X"FC82",X"FBF1",
		X"FC23",X"FA79",X"FC6A",X"FACD",X"FD22",X"FC2B",X"FD00",X"FC4C",X"FE0F",X"FE01",X"FE17",X"FEB4",X"FF2D",X"FFE6",X"FF13",X"010A",
		X"0053",X"0248",X"015F",X"02C7",X"0206",X"039A",X"0395",X"03A5",X"0359",X"050E",X"031B",X"059F",X"02AF",X"05A3",X"04E9",X"0534",
		X"0441",X"04DE",X"0530",X"0424",X"059F",X"03DC",X"06FA",X"036F",X"06E7",X"042C",X"06F8",X"0613",X"056E",X"057C",X"0411",X"0455",
		X"0354",X"02FF",X"0327",X"0246",X"02C7",X"0367",X"00CC",X"03EB",X"029F",X"03E8",X"0328",X"0160",X"03B1",X"02D9",X"00D6",X"03C2",
		X"001C",X"00F6",X"0170",X"FF6A",X"01D8",X"FFB2",X"0036",X"007F",X"FF6C",X"0023",X"006E",X"FE49",X"0297",X"FE3B",X"FEE8",X"02DE",
		X"FD62",X"0170",X"0137",X"FE63",X"00F2",X"FF82",X"FD73",X"FE67",X"FEB8",X"FCFA",X"FD6B",X"FE2E",X"FC4F",X"FDAE",X"FEF9",X"FD2A",
		X"FE2D",X"FE96",X"FE38",X"FEFE",X"FCCA",X"FEBD",X"FF1D",X"FC5F",X"FE0E",X"FE1E",X"FC14",X"FDB8",X"FF89",X"FDDD",X"FDD8",X"FF48",
		X"FF6C",X"FCCB",X"FFE2",X"0031",X"FC52",X"FF21",X"01BD",X"FD92",X"FD20",X"01EC",X"FF29",X"FD47",X"011D",X"01C4",X"FE3D",X"FFE2",
		X"03BD",X"FF5A",X"FFF9",X"034F",X"FF92",X"FF6C",X"0079",X"FF8C",X"FE5F",X"FEB8",X"FF44",X"FE56",X"FD0C",X"FFD0",X"0006",X"FD9F",
		X"FF37",X"0171",X"FF32",X"FE30",X"FFF9",X"0083",X"FEB8",X"FD08",X"0024",X"FF96",X"FBA9",X"FDA4",X"FFD0",X"FEBF",X"FB1C",X"FEFE",
		X"01E6",X"FD7B",X"FD98",X"02A2",X"027F",X"FC52",X"FEF3",X"036D",X"FE03",X"FB90",X"0201",X"00A8",X"FB04",X"FDCC",X"033C",X"FE4E",
		X"FB75",X"02F6",X"03BA",X"FC68",X"FF03",X"053C",X"0126",X"FBDF",X"0126",X"045E",X"FCC9",X"FC49",X"03B9",X"00AB",X"FAF4",X"FED6",
		X"03A0",X"FE28",X"FC3C",X"02B2",X"02FF",X"FCF9",X"FE9B",X"043F",X"00A2",X"FC50",X"0038",X"0498",X"FE00",X"FC4F",X"0222",X"0465",
		X"FE30",X"FDDF",X"049F",X"042F",X"FEBC",X"0045",X"049C",X"0191",X"FD9B",X"FF74",X"0104",X"FBED",X"FA1A",X"FE7F",X"FE1C",X"FB26",
		X"FC29",X"FECF",X"00D5",X"FFF8",X"01C0",X"02B3",X"02F3",X"03B9",X"051A",X"0381",X"0304",X"0519",X"0540",X"0385",X"0356",X"05A5",
		X"0671",X"05D3",X"0553",X"0704",X"06C1",X"0771",X"064D",X"04E6",X"055A",X"0750",X"05B7",X"0259",X"0409",X"0697",X"05C7",X"018D",
		X"0340",X"067B",X"054C",X"025C",X"033F",X"069E",X"04C4",X"02FB",X"0351",X"043E",X"0384",X"0253",X"0246",X"0178",X"0155",X"017B",
		X"0022",X"FEDD",X"FF9C",X"FFB9",X"FE4C",X"FD38",X"FD6A",X"FDA7",X"FBD4",X"FAF3",X"FB09",X"F9DF",X"F991",X"F8A3",X"F80D",X"F857",
		X"F7C8",X"F779",X"F795",X"F8A2",X"F89C",X"F87B",X"F84E",X"F84B",X"F9F9",X"F8F5",X"F783",X"F881",X"F9BF",X"F994",X"F6EA",X"F7CE",
		X"FAC9",X"F95B",X"F758",X"F911",X"FAEB",X"F9BC",X"F95C",X"FA68",X"FB01",X"FB9D",X"FC17",X"FC0D",X"FBEC",X"FC22",X"FD19",X"FC8D",
		X"FBA2",X"FCA2",X"FD3B",X"FD0D",X"FC63",X"FD05",X"FE43",X"FE83",X"FE46",X"FE5B",X"FFDC",X"FF35",X"FF1D",X"FF74",X"FFA5",X"FF88",
		X"FEBF",X"FF4B",X"FFBF",X"FE8A",X"FED7",X"00F7",X"00B1",X"0098",X"0152",X"02A2",X"02F8",X"02BA",X"02A7",X"0372",X"03DF",X"03A7",
		X"0311",X"0359",X"0528",X"04E7",X"0461",X"052C",X"06DD",X"0650",X"0542",X"0629",X"0772",X"0666",X"0597",X"06EE",X"0770",X"0666",
		X"0685",X"080C",X"0783",X"0711",X"0826",X"08CA",X"08A0",X"0867",X"09A5",X"09BA",X"090D",X"094B",X"09AB",X"09B1",X"0850",X"0836",
		X"08F5",X"0854",X"0754",X"075A",X"0802",X"0771",X"06A5",X"06A5",X"06DB",X"0674",X"05EC",X"058A",X"0450",X"0433",X"04C9",X"03A5",
		X"0202",X"01EC",X"02AA",X"0224",X"005E",X"0055",X"0176",X"009F",X"FEA3",X"FEDC",X"FF84",X"FED6",X"FDC9",X"FCEB",X"FCED",X"FC80",
		X"FB85",X"FB06",X"F9FF",X"F9D4",X"FA33",X"F90F",X"F8BA",X"F8DC",X"F90A",X"F8C0",X"F860",X"F8A0",X"F81B",X"F811",X"F747",X"F695",
		X"F5F2",X"F5BF",X"F58E",X"F4E1",X"F426",X"F46D",X"F591",X"F4D8",X"F421",X"F53B",X"F66E",X"F638",X"F52D",X"F685",X"F802",X"F656",
		X"F689",X"F76C",X"F7FA",X"F7AD",X"F778",X"F87F",X"F8D1",X"F928",X"FA15",X"FAC2",X"FA9C",X"FB4C",X"FBBA",X"FB4C",X"FBAD",X"FC60",
		X"FCE6",X"FBD6",X"FC3F",X"FDB3",X"FE58",X"FE4C",X"FEDB",X"001B",X"00D7",X"017E",X"01B3",X"027F",X"0303",X"0324",X"0382",X"0377",
		X"03A3",X"0381",X"03D3",X"0413",X"0409",X"04DB",X"0522",X"0520",X"056F",X"05DC",X"05EC",X"063F",X"0600",X"0682",X"062B",X"05B1",
		X"066A",X"0696",X"0702",X"0797",X"08DC",X"0985",X"0999",X"0AB6",X"0C8E",X"0CAB",X"0B7A",X"0BA5",X"0BF8",X"0AB5",X"0A04",X"0A1E",
		X"0989",X"07A2",X"069A",X"06BA",X"0650",X"060C",X"05BA",X"05AE",X"052C",X"0583",X"0530",X"0479",X"0489",X"0430",X"02F8",X"01D4",
		X"00BB",X"0104",X"011A",X"FFF0",X"FF73",X"FF25",X"FF60",X"FF7A",X"FEED",X"FEB4",X"FF8D",X"FFA3",X"FE1A",X"FDB0",X"FE00",X"FDE2",
		X"FD4A",X"FC6E",X"FCC7",X"FC95",X"FC54",X"FC82",X"FC77",X"FBEF",X"FC18",X"FB7D",X"FAED",X"FBE9",X"FC1A",X"FBDC",X"FB5A",X"FBFB",
		X"FB91",X"FBA3",X"FC04",X"FCCF",X"FCEF",X"FCC7",X"FD4A",X"FDD4",X"FE51",X"FE7A",X"FEB5",X"FE77",X"FE9C",X"FE6F",X"FF07",X"FEF3",
		X"FE93",X"FE88",X"FDEB",X"FDCE",X"FCE3",X"FC20",X"FC87",X"FC70",X"FB85",X"FBB0",X"FB73",X"FB4D",X"FBD2",X"FBBE",X"FBAA",X"FBD3",
		X"FC08",X"FB98",X"FB87",X"FB4D",X"FB56",X"FB71",X"FAD0",X"FA85",X"FAA9",X"FB86",X"FA34",X"FB42",X"FAF5",X"FBA4",X"FA7C",X"FBBE",
		X"FAD9",X"FB5B",X"FB87",X"FC9B",X"FC73",X"FCA5",X"FDB4",X"FDA1",X"FED3",X"FDB7",X"005B",X"FEC8",X"0110",X"FFF9",X"0214",X"0123",
		X"02CE",X"0266",X"02B3",X"0346",X"0474",X"024E",X"0458",X"035C",X"04F5",X"034D",X"04F9",X"04D3",X"0447",X"0577",X"0438",X"06DC",
		X"041C",X"0787",X"039D",X"073E",X"03E0",X"073D",X"058C",X"0520",X"0638",X"04F6",X"0646",X"045E",X"057A",X"0529",X"04BB",X"0458",
		X"0505",X"02F7",X"057A",X"02B8",X"03F3",X"036E",X"0232",X"0495",X"0204",X"0392",X"0524",X"01DC",X"03F2",X"0314",X"02E2",X"03B9",
		X"0063",X"0285",X"01B8",X"001B",X"015C",X"0102",X"0044",X"018A",X"FDF2",X"0173",X"00FB",X"FD83",X"02A4",X"FE8D",X"FEEA",X"0172",
		X"FDE5",X"FEC0",X"FFB9",X"FE37",X"FDE0",X"FEB1",X"FD51",X"FCDD",X"FE4C",X"FCF4",X"FBB4",X"FE29",X"FC55",X"FC26",X"FD99",X"FBB3",
		X"FDE8",X"FBE6",X"FB6E",X"FDD1",X"FB7A",X"FB42",X"FD9A",X"FBAD",X"FBB2",X"FDE5",X"FD06",X"FCC5",X"FE0A",X"0074",X"FDC7",X"FE2A",
		X"01EC",X"FF20",X"FCE4",X"0146",X"00B9",X"FBC9",X"FF96",X"0131",X"FD52",X"FD7C",X"0161",X"004D",X"FCC8",X"0142",X"0115",X"FD06",
		X"00DF",X"002A",X"FE0E",X"FF8B",X"FFAF",X"FEDD",X"FE4F",X"0011",X"0098",X"FE8F",X"FF19",X"01A6",X"FFA4",X"FE63",X"008D",X"0118",
		X"FEBA",X"FE9F",X"00DD",X"004B",X"FD7F",X"FECE",X"01D8",X"FEFA",X"FDB3",X"0067",X"028C",X"FEEC",X"FD6A",X"0305",X"023F",X"FD95",
		X"FF4E",X"03F2",X"FFA6",X"FC70",X"0145",X"01D5",X"FC26",X"FEB0",X"0310",X"FE15",X"FC10",X"0231",X"03B7",X"FC1A",X"FEA8",X"0500",
		X"0015",X"FC44",X"01D3",X"042A",X"FDB6",X"FC46",X"0305",X"01AC",X"FAD6",X"FF4D",X"03D6",X"FDED",X"FC78",X"0216",X"0271",X"FC5B",
		X"FE94",X"02E4",X"FF74",X"FB17",X"0057",X"027B",X"FC45",X"FB84",X"0161",X"01C6",X"FB5B",X"FDA2",X"0342",X"0266",X"FC75",X"0028",
		X"04BD",X"0167",X"FD29",X"003A",X"023C",X"FDC9",X"FBF9",X"FF72",X"FEE7",X"FA00",X"FC7E",X"0136",X"006D",X"FDEA",X"FF88",X"0369",
		X"0393",X"02ED",X"04E5",X"0431",X"032C",X"03CB",X"04E6",X"020A",X"0351",X"04BC",X"0429",X"02B6",X"03F6",X"069F",X"0725",X"06CC",
		X"0691",X"075C",X"0700",X"0843",X"072D",X"05B6",X"0675",X"0760",X"049B",X"0264",X"0562",X"07FF",X"062A",X"036C",X"0715",X"0937",
		X"0688",X"04DA",X"070C",X"078D",X"0438",X"0375",X"03AD",X"0336",X"01A6",X"0191",X"00E0",X"FEE5",X"FF33",X"FFD7",X"FE76",X"FE62",
		X"FF20",X"FEE3",X"FC9B",X"FB41",X"FC69",X"FBF1",X"FA2D",X"F917",X"F881",X"F87D",X"F74C",X"F618",X"F6E9",X"F787",X"F588",X"F595",
		X"F749",X"F785",X"F741",X"F7F3",X"F7C8",X"F86E",X"F899",X"F6F6",X"F6EA",X"F7B8",X"F93B",X"F742",X"F528",X"F744",X"F8B0",X"F684",
		X"F6A3",X"F911",X"F925",X"F88A",X"F90B",X"F9EE",X"F962",X"FA4B",X"FA99",X"F9D0",X"F8E4",X"F990",X"FAFA",X"FA73",X"FA58",X"FBE0",
		X"FD8F",X"FD76",X"FDA7",X"FEFD",X"003B",X"FFD9",X"FEEF",X"002D",X"001B",X"FEA1",X"FEEC",X"FF16",X"FEB7",X"FDA1",X"FE40",X"FEE4",
		X"FF36",X"FE62",X"011E",X"0234",X"0148",X"022F",X"0407",X"053C",X"0486",X"0467",X"04F2",X"064E",X"064A",X"0605",X"05B8",X"06E8",
		X"0702",X"06D4",X"0681",X"077D",X"08E7",X"07BD",X"070D",X"08A7",X"099D",X"07F1",X"0863",X"0A54",X"0A5E",X"093C",X"0A3A",X"0BC9",
		X"0A2C",X"0A2B",X"0B96",X"0BDC",X"0A1F",X"0A35",X"0B99",X"0A9E",X"0982",X"0A6A",X"0B32",X"099C",X"08C0",X"09C7",X"0A12",X"08F3",
		X"081D",X"08A4",X"0840",X"06CE",X"069C",X"069F",X"0597",X"0533",X"0502",X"04CF",X"0373",X"02E6",X"040B",X"02C1",X"0166",X"015F",
		X"0239",X"00A4",X"FEBE",X"FF2A",X"FFD9",X"FE5B",X"FCED",X"FDC9",X"FD86",X"FCF7",X"FC08",X"FC42",X"FB9C",X"FACB",X"FA78",X"F9FB",
		X"F85F",X"F82B",X"F82B",X"F6EE",X"F603",X"F5E2",X"F5F2",X"F507",X"F563",X"F53B",X"F501",X"F503",X"F57B",X"F57A",X"F4BD",X"F4A3",
		X"F516",X"F473",X"F351",X"F3F5",X"F543",X"F41F",X"F2D7",X"F3B9",X"F56A",X"F41F",X"F357",X"F5C4",X"F650",X"F5C0",X"F635",X"F777",
		X"F7E2",X"F79B",X"F842",X"F972",X"F950",X"F95C",X"FA6E",X"FABB",X"FA88",X"FB39",X"FC52",X"FB84",X"FBC3",X"FD40",X"FDB4",X"FDFC",
		X"FEC8",X"FFE3",X"FFE1",X"FFEC",X"00D8",X"01AF",X"0208",X"0287",X"026D",X"0337",X"043E",X"03EF",X"040D",X"0487",X"04C3",X"0479",
		X"04FE",X"053B",X"0547",X"04FA",X"0544",X"05A7",X"061E",X"05DF",X"063E",X"0712",X"0734",X"07AD",X"0726",X"07E6",X"0872",X"08DB",
		X"094F",X"0A6B",X"0AB9",X"0B24",X"0B70",X"0CF3",X"0DFA",X"0CFB",X"0C1E",X"0CAA",X"0CBE",X"0B51",X"0A62",X"0986",X"08B0",X"0766",
		X"0771",X"068C",X"0610",X"05F1",X"05FC",X"0471",X"0484",X"05BF",X"0423",X"02D0",X"0268",X"02EB",X"022C",X"FFF2",X"FFFD",X"FFD8",
		X"FE43",X"FE75",X"FE65",X"FDCB",X"FEA1",X"FED4",X"FDDA",X"FD6A",X"FEDF",X"FEA4",X"FDBC",X"FD98",X"FD71",X"FC9C",X"FBB2",X"FB0E",
		X"FB3E",X"FA97",X"F98B",X"F934",X"F8D7",X"F878",X"F8E3",X"F92E",X"F94A",X"F9C2",X"F9D6",X"FA04",X"F9FB",X"FA58",X"FAF7",X"FAF8",
		X"FAF9",X"FAF8",X"FB67",X"FBFC",X"FC65",X"FD40",X"FCF3",X"FD1C",X"FDF6",X"FDCE",X"FDF7",X"FE16",X"FEA5",X"FE6F",X"FDC4",X"FD8F",
		X"FD43",X"FD4B",X"FC6C",X"FC22",X"FC53",X"FC20",X"FBC5",X"FB9C",X"FC10",X"FC6D",X"FCA3",X"FCAF",X"FCFC",X"FDAE",X"FDD5",X"FD90",
		X"FD75",X"FD49",X"FDDC",X"FD2C",X"FD2F",X"FCD4",X"FD16",X"FD7C",X"FD30",X"FD5A",X"FD0C",X"FDCE",X"FDA4",X"FF3F",X"FD07",X"FF12",
		X"FE82",X"0082",X"FEF2",X"0039",X"002A",X"01B0",X"00B1",X"01CE",X"0277",X"032E",X"03F5",X"0314",X"049A",X"040C",X"0597",X"0522",
		X"04FA",X"0567",X"05F5",X"046E",X"061F",X"03E2",X"076E",X"041E",X"06A7",X"0490",X"06CC",X"051A",X"06B7",X"0614",X"07B0",X"07BC",
		X"05BD",X"0856",X"052A",X"087C",X"0476",X"0685",X"04F1",X"0520",X"04BC",X"03B6",X"035C",X"042E",X"026C",X"0348",X"0231",X"01AD",
		X"036D",X"00B2",X"02F6",X"01B9",X"0184",X"0305",X"0024",X"011E",X"01DB",X"FEF4",X"0183",X"FE08",X"FEF2",X"FF35",X"FCE6",X"FE8D",
		X"FD68",X"FCF0",X"FE5B",X"FCE7",X"FD3C",X"FF5A",X"FABE",X"FF8A",X"FD10",X"FA8B",X"FFC6",X"FAF8",X"FBC4",X"FDA1",X"FB79",X"FBB1",
		X"FD0D",X"FC44",X"FB68",X"FD6F",X"FC81",X"FBC3",X"FD0F",X"FBF3",X"FA4C",X"FC52",X"FAF4",X"FB59",X"FB36",X"F9DD",X"FC87",X"FABB",
		X"FADB",X"FDF8",X"FC8E",X"FC49",X"FEA5",X"FDBE",X"FDA5",X"FF14",X"FFBD",X"FE52",X"FE37",X"0132",X"FF1C",X"FE5B",X"01A9",X"0002",
		X"FD81",X"0201",X"01E4",X"FE81",X"0189",X"039A",X"0107",X"FF0F",X"03E2",X"02B7",X"FDCA",X"0239",X"0258",X"FE70",X"009A",X"0079",
		X"005A",X"0085",X"0167",X"0189",X"0033",X"01A7",X"027F",X"0046",X"FFDB",X"02B7",X"010C",X"FEAA",X"FFAB",X"0210",X"00F2",X"FF01",
		X"0127",X"0395",X"005B",X"FFD3",X"0321",X"0288",X"0050",X"FFB2",X"0449",X"00BA",X"FD75",X"009A",X"0360",X"FE32",X"FC81",X"034B",
		X"0173",X"FBF8",X"FFC6",X"038D",X"FD7D",X"FCB4",X"028A",X"01B5",X"FB5C",X"FFF2",X"042E",X"FE09",X"FCB5",X"0355",X"0316",X"FCD1",
		X"FED8",X"04BF",X"00D8",X"FC2F",X"019F",X"037A",X"FC61",X"FD31",X"031A",X"002F",X"FBAC",X"0083",X"02D4",X"FE29",X"FD33",X"0339",
		X"0292",X"FCE1",X"FF5E",X"0451",X"0103",X"FCD7",X"0130",X"0498",X"FEF7",X"FC30",X"01C0",X"03FA",X"FE18",X"FD92",X"03A5",X"0326",
		X"FE73",X"FEAD",X"029D",X"FF8D",X"FC49",X"FEFA",X"FFEF",X"FB38",X"FABB",X"FE5C",X"003B",X"FD2A",X"FCA3",X"FFAA",X"00A2",X"0115",
		X"02C4",X"0212",X"0046",X"0260",X"03DB",X"0191",X"00C8",X"03D1",X"0366",X"01F4",X"01DA",X"0482",X"04DF",X"04CF",X"05E0",X"0425",
		X"041A",X"0681",X"06D0",X"042E",X"0414",X"063D",X"05A1",X"0164",X"0119",X"0543",X"051F",X"01E5",X"021D",X"0447",X"0450",X"01F6",
		X"02AE",X"0403",X"0352",X"018C",X"019F",X"022F",X"00C8",X"01E5",X"0104",X"FF52",X"FEB0",X"FFDF",X"FE59",X"FD16",X"FDF9",X"FEC1",
		X"FC7B",X"FA76",X"FC70",X"FC4B",X"FB0E",X"FA89",X"FA73",X"F9DC",X"F935",X"F869",X"F8FB",X"F919",X"F8BF",X"F836",X"F811",X"F87C",
		X"F9B9",X"FA32",X"F8C8",X"F902",X"FACB",X"F9D5",X"F815",X"F7F1",X"FB51",X"FA28",X"F70B",X"F7CC",X"FA43",X"F973",X"F7E4",X"F995",
		X"FA7D",X"FADE",X"FB2D",X"FACD",X"FAC6",X"FBD0",X"FCCB",X"FCEA",X"FB93",X"FC6A",X"FD39",X"FD7F",X"FD34",X"FD7C",X"FF08",X"FF27",
		X"FEBA",X"FECA",X"004A",X"00B9",X"FFCA",X"0065",X"00F8",X"00A2",X"FFFE",X"00FE",X"019A",X"003A",X"FFCE",X"0142",X"017A",X"0024",
		X"0110",X"022E",X"028D",X"0230",X"02E0",X"0428",X"0500",X"0495",X"0485",X"0528",X"069F",X"0692",X"0605",X"0681",X"0777",X"07D5",
		X"0689",X"067C",X"0799",X"0796",X"0669",X"0679",X"070E",X"063A",X"057C",X"073A",X"082D",X"06D9",X"073E",X"089E",X"0817",X"0808",
		X"08F9",X"09CE",X"0825",X"06B1",X"081F",X"0839",X"0745",X"0665",X"0761",X"06D3",X"05A2",X"0604",X"06E3",X"06E6",X"0587",X"0663",
		X"061E",X"055E",X"04A8",X"04A9",X"0409",X"0333",X"035A",X"02EF",X"0167",X"005D",X"015A",X"00F5",X"FE83",X"FE06",X"FEF8",X"FEAE",
		X"FC78",X"FC9D",X"FDFE",X"FD72",X"FC53",X"FC5A",X"FC2D",X"FCAD",X"FBE6",X"FB51",X"FB05",X"FA97",X"FA8B",X"FA74",X"F93D",X"F962",
		X"FA92",X"F9CE",X"F8F1",X"F91C",X"F87E",X"F87E",X"F814",X"F71C",X"F724",X"F630",X"F68E",X"F608",X"F5CC",X"F5E8",X"F73D",X"F6EA",
		X"F63C",X"F6D1",X"F8A9",X"F88E",X"F724",X"F807",X"F97C",X"F85C",X"F6FC",X"F8C9",X"F8F8",X"F83B",X"F88B",X"F968",X"F9AF",X"FA4A",
		X"FAC4",X"FB77",X"FC57",X"FC8E",X"FD91",X"FD3E",X"FD00",X"FE02",X"FEC6",X"FE27",X"FD60",X"FE56",X"FF09",X"FE88",X"FE9C",X"FFFF",
		X"003E",X"0026",X"00F7",X"022B",X"02DA",X"02F5",X"0348",X"03B6",X"035D",X"0349",X"03D7",X"037A",X"0327",X"0331",X"03A5",X"0398",
		X"0496",X"05AC",X"05FF",X"0638",X"0711",X"0744",X"07B1",X"0798",X"07F7",X"088B",X"07F0",X"07CD",X"086B",X"0961",X"0925",X"0970",
		X"0AF0",X"0BD6",X"0AAC",X"0B7D",X"0C38",X"0AD8",X"0987",X"09EC",X"0957",X"074B",X"05A1",X"05C7",X"0566",X"04E4",X"042D",X"02FC",
		X"0251",X"0222",X"022B",X"019D",X"0192",X"017B",X"0103",X"FFF1",X"FFD4",X"FFE6",X"FFE8",X"FEC8",X"FE94",X"FE8A",X"FE05",X"FDDC",
		X"FDB9",X"FD30",X"FDB8",X"FE7F",X"FD49",X"FC73",X"FD43",X"FE10",X"FDDB",X"FD17",X"FCCD",X"FD0C",X"FBFC",X"FB87",X"FBD7",X"FBA5",
		X"FA59",X"FA32",X"FA01",X"F9BA",X"FA2C",X"FB12",X"FB05",X"FB74",X"FC28",X"FC5E",X"FCAA",X"FD38",X"FEBE",X"FEAF",X"FE65",X"FED2",
		X"FFAD",X"FEF3",X"FFA3",X"0058",X"FF8A",X"FEF2",X"FF5A",X"001A",X"FFAE",X"FFC9",X"0085",X"0024",X"FF65",X"FE7C",X"FE6E",X"FECD",
		X"FE12",X"FD67",X"FD2D",X"FCEB",X"FCB2",X"FCFA",X"FD3C",X"FDA1",X"FD23",X"FCBE",X"FD13",X"FD26",X"FCBB",X"FCFB",X"FCFC",X"FC34",
		X"FB9D",X"FB9B",X"FBAA",X"FADD",X"FBE6",X"FB98",X"FBD1",X"FB4A",X"FCD5",X"FB76",X"FD3E",X"FD2D",X"FD90",X"FC0B",X"FDA3",X"FD81",
		X"FD66",X"FD7E",X"FDCC",X"FE8D",X"FDBE",X"FF90",X"FF2C",X"0108",X"0094",X"023B",X"01AE",X"0270",X"02D8",X"03B1",X"0298",X"0478",
		X"0254",X"04FE",X"0222",X"04DB",X"0305",X"048B",X"02EC",X"043E",X"045D",X"0407",X"056B",X"03BE",X"0763",X"0391",X"072C",X"039E",
		X"06D8",X"04D5",X"056C",X"04E8",X"0381",X"04F4",X"03C2",X"0302",X"045D",X"035E",X"0389",X"044E",X"0236",X"0483",X"02AF",X"03A9",
		X"0333",X"00C3",X"0302",X"0120",X"001B",X"0278",X"FFBC",X"0149",X"0043",X"FFB5",X"01C4",X"FFF4",X"008D",X"00EC",X"001B",X"0139",
		X"0041",X"FE8E",X"031F",X"FDEB",X"FE87",X"01C2",X"FBD9",X"005B",X"FEC0",X"FCA1",X"FF7C",X"FE57",X"FD6B",X"FE66",X"FEF6",X"FD45",
		X"FE18",X"FED4",X"FC87",X"FD78",X"FEB5",X"FBF4",X"FDC6",X"FD67",X"FC19",X"FDBE",X"FBEA",X"FDF6",X"FD93",X"FB78",X"FE2D",X"FE2A",
		X"FC59",X"FEBE",X"FF8A",X"FD6B",X"FE35",X"0014",X"FFE6",X"FD32",X"0176",X"01BF",X"FD88",X"000E",X"0347",X"FF32",X"FEAA",X"0301",
		X"0071",X"FDF0",X"013A",X"027B",X"FE36",X"FFC6",X"0312",X"FE13",X"FF07",X"0325",X"FF1C",X"FFE1",X"0150",X"00CD",X"0053",X"0130",
		X"01E9",X"00B6",X"FF95",X"01E4",X"0196",X"FECF",X"003F",X"01C5",X"0014",X"FECE",X"012D",X"01B1",X"FF86",X"FF19",X"023A",X"017D",
		X"FE51",X"0049",X"0278",X"00B5",X"FD18",X"00B7",X"02E4",X"FE0B",X"FD4B",X"01A3",X"016D",X"FC5F",X"FEFC",X"02D4",X"FE4F",X"FC1A",
		X"0223",X"0054",X"FB73",X"FF06",X"02FC",X"FD53",X"FAEA",X"022E",X"018D",X"FAF4",X"FE95",X"0379",X"FF5B",X"FBF0",X"00D1",X"030B",
		X"FC9A",X"FC47",X"0232",X"FF48",X"FA04",X"FE82",X"01FB",X"FCC0",X"FBB4",X"01C7",X"014B",X"FC8B",X"FE57",X"03DB",X"FFB8",X"FC27",
		X"004C",X"0304",X"FDB8",X"FB5C",X"0186",X"02C4",X"FC7E",X"FC74",X"0351",X"0213",X"FCAA",X"FEA7",X"0338",X"0046",X"FC4C",X"FEAE",
		X"00F1",X"FCDB",X"FB43",X"0004",X"FFB2",X"FCD3",X"FD65",X"009F",X"01D5",X"0017",X"01DF",X"02B7",X"0270",X"03AB",X"0528",X"03B3",
		X"039E",X"0613",X"05BA",X"046B",X"04A9",X"068D",X"0698",X"0639",X"0577",X"0615",X"0620",X"0693",X"058C",X"0428",X"05A1",X"0676",
		X"04F8",X"01FB",X"0419",X"06F4",X"05C7",X"025B",X"0478",X"07BD",X"060E",X"03BD",X"0523",X"070E",X"04E1",X"034F",X"0437",X"04CD",
		X"03C9",X"02C3",X"02FA",X"0222",X"020D",X"0289",X"00DB",X"0051",X"0070",X"0016",X"FE76",X"FDDA",X"FD8C",X"FD02",X"FAE4",X"FA96",
		X"FA9C",X"FA58",X"F9E2",X"F8F0",X"F943",X"F9A5",X"F922",X"F804",X"F891",X"F885",X"F7FF",X"F7C0",X"F74B",X"F73A",X"F815",X"F7B2",
		X"F6A0",X"F864",X"F92F",X"F855",X"F717",X"F7EC",X"FAB4",X"F892",X"F6F2",X"F857",X"F92F",X"F81F",X"F7C6",X"F80F",X"F84E",X"F8A3",
		X"F98D",X"F948",X"F8F6",X"F9B6",X"FB17",X"FAF3",X"FA55",X"FB51",X"FC70",X"FC65",X"FBDF",X"FBDD",X"FCCA",X"FD5F",X"FC86",X"FC40",
		X"FDD0",X"FD10",X"FC6F",X"FD5E",X"FDAF",X"FD53",X"FD29",X"FE54",X"FE6F",X"FE11",X"FF18",X"0164",X"0048",X"011A",X"0220",X"02FA",
		X"039E",X"033D",X"0457",X"0548",X"05C4",X"056D",X"0529",X"05E1",X"072B",X"064F",X"05BD",X"0687",X"079B",X"06D8",X"05F3",X"0728",
		X"08BA",X"0779",X"06F7",X"08CC",X"09E3",X"08F2",X"0890",X"0A81",X"09AF",X"0979",X"0AA2",X"0B5F",X"0AA7",X"0A54",X"0B20",X"0B1F",
		X"09F4",X"0A70",X"0AFE",X"0A29",X"08CE",X"0935",X"0A49",X"0992",X"08E6",X"0931",X"09B1",X"088B",X"0812",X"083D",X"081D",X"07C8",
		X"0744",X"05A3",X"04BB",X"040B",X"0495",X"0329",X"0165",X"0138",X"021A",X"017D",X"FFB0",X"002B",X"015A",X"009F",X"FEC2",X"FF3C",
		X"FFD3",X"FF17",X"FE0C",X"FE07",X"FE0C",X"FD33",X"FC91",X"FC50",X"FB6F",X"FAB3",X"FAF2",X"F9E0",X"F8C6",X"F8DC",X"F938",X"F894",
		X"F78F",X"F790",X"F71F",X"F6A3",X"F630",X"F636",X"F565",X"F4EE",X"F54A",X"F4C8",X"F44C",X"F475",X"F55B",X"F503",X"F41D",X"F518",
		X"F582",X"F528",X"F3D8",X"F4EC",X"F601",X"F472",X"F419",X"F4C5",X"F57D",X"F53A",X"F54C",X"F660",X"F6FB",X"F71F",X"F742",X"F838",
		X"F8A5",X"F98C",X"F9C5",X"F9B9",X"F9E9",X"FA40",X"FB70",X"FA56",X"FAE3",X"FC26",X"FCD6",X"FD34",X"FD79",X"FE50",X"FF82",X"008D",
		X"0104",X"019C",X"0223",X"0271",X"0294",X"02EC",X"0369",X"035A",X"038D",X"03E5",X"0402",X"0477",X"0504",X"0571",X"060C",X"067B",
		X"06AC",X"0712",X"074F",X"07BA",X"07AE",X"0797",X"082A",X"087E",X"087B",X"08F3",X"0A2B",X"0A95",X"0ACD",X"0BBB",X"0D47",X"0D3F",
		X"0C95",X"0D0A",X"0D27",X"0C12",X"0BA5",X"0B43",X"0A52",X"0943",X"0858",X"0813",X"07C4",X"0799",X"074D",X"0709",X"0677",X"0706",
		X"06C3",X"05A9",X"054C",X"055C",X"0499",X"02E5",X"01CD",X"01FF",X"01D0",X"0082",X"000A",X"0027",X"0074",X"0088",X"0035",X"FFEE",
		X"0003",X"0058",X"FF0B",X"FE8E",X"FE1A",X"FDE5",X"FCDB",X"FBDF",X"FB8B",X"FB14",X"FAA5",X"FAA9",X"FA8F",X"FA55",X"FAF6",X"FAC8",
		X"FA86",X"FB09",X"FB91",X"FB97",X"FB63",X"FB6F",X"FBAB",X"FBAA",X"FBD0",X"FC6B",X"FC8B",X"FC19",X"FC69",X"FC4D",X"FCCF",X"FD41",
		X"FD5F",X"FD78",X"FD1E",X"FCE5",X"FD12",X"FD03",X"FC68",X"FC6B",X"FBBE",X"FB93",X"FA3F",X"F9AB",X"F9FE",X"F9DD",X"F989",X"F9B0",
		X"FA02",X"FA4F",X"FAB9",X"FA9E",X"FB5F",X"FB08",X"FB50",X"FADF",X"FA86",X"FA4E",X"FA53",X"FAFB",X"FA83",X"FA35",X"FA27",X"FB2F",
		X"FA00",X"FAED",X"FA5F",X"FBB9",X"FA64",X"FB6F",X"FB18",X"FBD5",X"FC0C",X"FCA3",X"FCC1",X"FCC6",X"FE99",X"FE9B",X"FF69",X"FE54",
		X"01A9",X"006C",X"0290",X"015C",X"0419",X"0340",X"0444",X"0464",X"04CC",X"04C7",X"05C5",X"03DF",X"05D3",X"0413",X"0596",X"042A",
		X"0502",X"0594",X"054F",X"06B3",X"0518",X"084D",X"0657",X"096F",X"0558",X"09CA",X"06F2",X"08EE",X"06ED",X"06EA",X"07B1",X"066F",
		X"07F4",X"056A",X"06D8",X"0602",X"068B",X"05ED",X"066A",X"053F",X"074D",X"0516",X"0579",X"0579",X"03C2",X"064F",X"028F",X"02FB",
		X"043D",X"017E",X"02EB",X"01B7",X"0076",X"028E",X"FF81",X"0131",X"0048",X"FF26",X"00D1",X"FF91",X"FFD3",X"0172",X"FE97",X"0094",
		X"00DD",X"FDAF",X"02FC",X"FE76",X"FE00",X"00C0",X"FDE0",X"FE73",X"FE97",X"FD56",X"FCF1",X"FDAB",X"FC54",X"FBC2",X"FD71",X"FC0D",
		X"FA6D",X"FC19",X"FACD",X"FA07",X"FB96",X"F9F9",X"FB6E",X"FA80",X"FA22",X"FCA0",X"FAF4",X"FB69",X"FDB8",X"FC89",X"FB6F",X"FE66",
		X"FDD7",X"FBDC",X"FD53",X"FEBF",X"FC4A",X"FB57",X"FF4D",X"FD51",X"FAEC",X"FFC9",X"0045",X"FB94",X"FF6B",X"0116",X"FDE6",X"FE8D",
		X"01AD",X"FFED",X"FCAA",X"00D3",X"FFE2",X"FB93",X"FF3A",X"FEDD",X"FCC3",X"FE54",X"FEF4",X"FE0C",X"FD42",X"FFA0",X"0026",X"FE3E",
		X"FED8",X"022D",X"FFB9",X"FE78",X"0074",X"013D",X"FEF2",X"FEC9",X"0142",X"0100",X"FE74",X"FF1F",X"02B3",X"0005",X"FEED",X"0118",
		X"038B",X"FF97",X"FD62",X"0304",X"027B",X"FD2A",X"FE9F",X"0369",X"FFD5",X"FC93",X"0206",X"03CE",X"FD79",X"FFFC",X"04B1",X"007F",
		X"FCDD",X"02C5",X"0482",X"FD12",X"FECA",X"05C0",X"0102",X"FC6F",X"023E",X"0560",X"FF4A",X"FE27",X"04D2",X"0357",X"FCC6",X"0074",
		X"0521",X"FFDA",X"FD3D",X"02CE",X"0399",X"FD33",X"FF38",X"0482",X"025B",X"FCD0",X"019A",X"0438",X"FF58",X"FD84",X"03C1",X"03FE",
		X"FD00",X"FEAB",X"04AC",X"031C",X"FC9B",X"0099",X"04D1",X"0142",X"FCFF",X"00B5",X"01CE",X"FDEB",X"FBCA",X"FF63",X"FF03",X"FA3C",
		X"FBE3",X"00B9",X"003F",X"FCF4",X"FE63",X"0209",X"0243",X"00FC",X"032B",X"025A",X"0234",X"02F3",X"03DD",X"0174",X"030E",X"046C",
		X"038B",X"01C3",X"02C8",X"0499",X"04F3",X"0465",X"03E5",X"0435",X"0373",X"0565",X"042A",X"02B3",X"04A5",X"067C",X"0390",X"013E",
		X"0481",X"07C2",X"04DA",X"0189",X"04A2",X"066F",X"03E8",X"022D",X"0422",X"0518",X"0227",X"0177",X"01CE",X"0247",X"01C9",X"019D",
		X"00DC",X"FFAB",X"FFD1",X"001C",X"FDE1",X"FD54",X"FDF1",X"FD90",X"FAF3",X"F9C7",X"FB55",X"FAF4",X"F941",X"F909",X"F911",X"F8CB",
		X"F8A8",X"F822",X"F8FD",X"F905",X"F772",X"F73D",X"F7D0",X"F7CC",X"F789",X"F7F3",X"F86D",X"F8A6",X"F96B",X"F835",X"F7EA",X"F938",
		X"FAD8",X"F8E0",X"F72B",X"F9B8",X"FAF7",X"F897",X"F82D",X"FA2E",X"FA11",X"F942",X"F9C8",X"FA62",X"F9CC",X"FB10",X"FC00",X"FB22",
		X"FA7F",X"FBC2",X"FCCF",X"FBFD",X"FBF0",X"FD9E",X"FE4D",X"FDEE",X"FE09",X"FF33",X"0064",X"0016",X"FF05",X"0090",X"0105",X"000C",
		X"0083",X"011D",X"0110",X"002A",X"0105",X"022B",X"01E3",X"00CF",X"0356",X"03BC",X"0243",X"02E9",X"0473",X"051E",X"0463",X"0466",
		X"054D",X"06BF",X"0779",X"06FC",X"06FF",X"086E",X"08A9",X"07AF",X"078E",X"0889",X"0944",X"07E0",X"06A5",X"07A5",X"08C5",X"0760",
		X"06EC",X"091A",X"0A37",X"0881",X"0904",X"0B0F",X"0AA1",X"0ACA",X"0B10",X"0B60",X"0987",X"0970",X"0A39",X"0876",X"0783",X"073E",
		X"0761",X"063C",X"052F",X"067E",X"06C1",X"05D3",X"053D",X"0638",X"062D",X"0517",X"03A7",X"036B",X"032F",X"02CB",X"01F4",X"00C0",
		X"00B1",X"00A3",X"0114",X"FFF4",X"FF40",X"FF9B",X"00D8",X"FFE1",X"FE1A",X"FE69",X"FF79",X"FDA9",X"FBBF",X"FC7A",X"FCB4",X"FB3E",
		X"FA49",X"FAA6",X"FAC6",X"F9FD",X"F970",X"F92F",X"F88D",X"F8A6",X"F916",X"F80D",X"F714",X"F71A",X"F6C9",X"F648",X"F5E4",X"F554",
		X"F4F0",X"F49C",X"F53D",X"F4AF",X"F474",X"F55C",X"F612",X"F606",X"F5B0",X"F6C5",X"F768",X"F6D0",X"F5C2",X"F642",X"F736",X"F6B6",
		X"F57C",X"F79F",X"F7D9",X"F6E5",X"F77B",X"F8E7",X"F96A",X"F933",X"FA62",X"FB16",X"FB14",X"FAAD",X"FBB3",X"FB84",X"FB4E",X"FC9E",
		X"FCCD",X"FC31",X"FC9C",X"FEAB",X"FF0B",X"FF18",X"0036",X"0101",X"012B",X"0159",X"023B",X"02E6",X"033D",X"0348",X"02F3",X"032E",
		X"034F",X"0447",X"0434",X"03EF",X"045D",X"042C",X"04A0",X"0546",X"05FE",X"05FF",X"0667",X"06CC",X"0770",X"0702",X"079A",X"07D6",
		X"07C6",X"0813",X"07D5",X"0891",X"08EB",X"093B",X"0A99",X"0B3B",X"0B66",X"0C54",X"0CD8",X"0D68",X"0DD3",X"0CE9",X"0BBE",X"0B97",
		X"0B5B",X"095D",X"083B",X"0800",X"06F4",X"061D",X"0601",X"05DE",X"054F",X"0571",X"0567",X"04AE",X"040B",X"0473",X"03B1",X"0227",
		X"012C",X"0109",X"0080",X"FEAB",X"FEDE",X"FF25",X"FE8E",X"FE29",X"FD5E",X"FE15",X"FE39",X"FEF8",X"FDA8",X"FC89",X"FD4C",X"FD42",
		X"FC5F",X"FBCD",X"FBB3",X"FB92",X"FB21",X"FA3C",X"FB3A",X"FB19",X"FAAD",X"FA7D",X"FA18",X"FAAD",X"FA7B",X"FA76",X"FAFB",X"FAC1",
		X"FAB2",X"FA9E",X"FAE7",X"FB6E",X"FBE7",X"FBF5",X"FC05",X"FC56",X"FD0A",X"FD3E",X"FD02",X"FD73",X"FD1F",X"FD25",X"FCE0",X"FCC4",
		X"FD15",X"FCCF",X"FD6D",X"FC9D",X"FC76",X"FC0F",X"FBBA",X"FBE9",X"FBF5",X"FBAB",X"FC06",X"FC1D",X"FC0C",X"FC27",X"FBF4",X"FC77",
		X"FC13",X"FC4E",X"FCA9",X"FC96",X"FC6E",X"FC54",X"FC54",X"FB88",X"FCF5",X"FCC9",X"FC72",X"FBA6",X"FCA0",X"FD63",X"FCC3",X"FCEC",
		X"FDB1",X"FE0E",X"FD4E",X"FEB1",X"FD86",X"FF42",X"FE45",X"0047",X"FE45",X"0008",X"FF7F",X"0125",X"0003",X"0136",X"01BB",X"0274",
		X"02E9",X"0307",X"046F",X"0439",X"059A",X"055D",X"0535",X"05DD",X"0550",X"0432",X"05CF",X"037E",X"05FD",X"036A",X"05CD",X"0372",
		X"0669",X"0409",X"06A8",X"050A",X"06D1",X"066E",X"05A9",X"0783",X"049E",X"0877",X"04BC",X"073C",X"056B",X"0676",X"04EE",X"0461",
		X"04F4",X"04CC",X"0307",X"03D6",X"02A8",X"0233",X"0300",X"00C9",X"037E",X"00D4",X"00DD",X"026C",X"FF72",X"0107",X"00C6",X"FE49",
		X"010D",X"FE48",X"0001",X"FF26",X"FDCE",X"0002",X"FF28",X"FE80",X"FFEE",X"FE2B",X"FF40",X"002E",X"FBA6",X"0185",X"FDCB",X"FCCE",
		X"0141",X"FD20",X"FE9E",X"FF46",X"FD1D",X"FD57",X"FE73",X"FD2E",X"FBE7",X"FD6F",X"FC1C",X"FAB3",X"FC2C",X"FB2E",X"FA3E",X"FC62",
		X"FAA1",X"FC4A",X"FB16",X"FAC5",X"FD89",X"FB2E",X"FC53",X"FE89",X"FD32",X"FD2E",X"FEC5",X"FE2A",X"FE74",X"0013",X"FFF5",X"FE74",
		X"FF13",X"0191",X"FE19",X"FE24",X"0224",X"FF02",X"FD1B",X"00F6",X"009C",X"FCF9",X"006E",X"01A5",X"FEC7",X"FDD8",X"02F3",X"014C",
		X"FD2A",X"0335",X"0199",X"FF04",X"0299",X"01ED",X"00AA",X"0050",X"0158",X"0129",X"FFAA",X"0021",X"01A3",X"FE54",X"FEDD",X"0143",
		X"0029",X"FEBF",X"0000",X"01B0",X"0045",X"FF20",X"00C1",X"01FD",X"FE96",X"FF87",X"01AD",X"0074",X"FE5E",X"FEE3",X"0323",X"FF92",
		X"FD1E",X"00D1",X"02A7",X"FE1B",X"FDBC",X"0363",X"00DF",X"FC09",X"00C6",X"028A",X"FC67",X"FD41",X"0224",X"FFF4",X"FA42",X"0043",
		X"032A",X"FC90",X"FD1D",X"0363",X"0161",X"FBA4",X"FFB6",X"04C6",X"FF4D",X"FC7B",X"0269",X"02BA",X"FBCE",X"FE3E",X"0380",X"FF42",
		X"FB3C",X"0101",X"0203",X"FCD1",X"FDEE",X"044A",X"0253",X"FCDB",X"00AB",X"0517",X"0075",X"FD45",X"0273",X"03ED",X"FE18",X"FC74",
		X"01E5",X"035A",X"FDB1",X"FE93",X"03B3",X"02A9",X"FE22",X"FF93",X"02A0",X"FEE1",X"FBAE",X"FECE",X"FE8B",X"F9D2",X"FAC1",X"FE8C",
		X"0052",X"FD23",X"FE71",X"0106",X"0178",X"0305",X"0548",X"02BC",X"0184",X"03E3",X"048F",X"0272",X"02A2",X"059F",X"0441",X"02B5",
		X"033F",X"05FE",X"0691",X"0661",X"06B2",X"0563",X"0560",X"0873",X"07C2",X"04C6",X"063F",X"08EE",X"07BC",X"0344",X"04F6",X"0930",
		X"0841",X"03A7",X"04C1",X"0707",X"05B9",X"02C0",X"03D5",X"04DC",X"02FF",X"01C8",X"023A",X"0267",X"017F",X"02C2",X"020F",X"0049",
		X"0030",X"0150",X"FF3E",X"FE79",X"FEDE",X"FF58",X"FCCD",X"FAFD",X"FC5B",X"FC0E",X"FB44",X"FA71",X"F9F6",X"F98F",X"F957",X"F903",
		X"F94C",X"F8F7",X"F824",X"F83B",X"F741",X"F6FA",X"F822",X"F8CB",X"F754",X"F858",X"F9E5",X"F8B8",X"F713",X"F770",X"FA9E",X"F8D0",
		X"F615",X"F755",X"F8DA",X"F766",X"F689",X"F766",X"F7A9",X"F798",X"F879",X"F810",X"F7AF",X"F9AD",X"FB02",X"FB40",X"FA46",X"FAF1",
		X"FCC4",X"FC55",X"FBF3",X"FC68",X"FD1A",X"FD51",X"FC8A",X"FCA1",X"FD9D",X"FD60",X"FC68",X"FD97",X"FDD5",X"FD29",X"FD31",X"FE10",
		X"FE8C",X"FDB3",X"FDC0",X"FFC6",X"FF9C",X"FE53",X"FFD8",X"00BB",X"0138",X"00B8",X"0205",X"0385",X"0468",X"03AE",X"03BA",X"04CF",
		X"0617",X"0631",X"0505",X"057E",X"06B8",X"0615",X"04ED",X"0585",X"06BF",X"0608",X"04D3",X"05E3",X"0780",X"0693",X"062D",X"0884",
		X"09F0",X"08DE",X"0995",X"0AF9",X"0ABF",X"0A70",X"0BCA",X"0C41",X"0ACD",X"0B3D",X"0AF5",X"0A7B",X"0A35",X"0A1D",X"0ACF",X"09D7",
		X"08D1",X"09CC",X"0A1F",X"09A1",X"08B3",X"08C2",X"08F6",X"085E",X"0745",X"06B1",X"0576",X"0502",X"0560",X"04B8",X"0369",X"03C3",
		X"0422",X"0397",X"01F1",X"025A",X"0378",X"0328",X"010A",X"0148",X"021B",X"008E",X"FF84",X"FF1C",X"FE5A",X"FE2E",X"FD3A",X"FC49",
		X"FC0D",X"FB74",X"FB9B",X"FB83",X"FABB",X"FACB",X"FAC1",X"F9FE",X"F9B9",X"F91C",X"F896",X"F85F",X"F78E",X"F652",X"F570",X"F53C",
		X"F5B0",X"F4DE",X"F453",X"F3F6",X"F52D",X"F451",X"F379",X"F4AE",X"F5B2",X"F501",X"F420",X"F4AA",X"F5D0",X"F4FF",X"F408",X"F5A2",
		X"F55F",X"F512",X"F614",X"F6AC",X"F6CD",X"F769",X"F7E9",X"F83B",X"F859",X"F86F",X"F93D",X"F89C",X"F8B9",X"FA00",X"F9A2",X"F952",
		X"F8ED",X"FADA",X"FB23",X"FB83",X"FC79",X"FD50",X"FE04",X"FEDC",X"FFB0",X"006C",X"0200",X"016A",X"0199",X"0123",X"01B8",X"022B",
		X"018A",X"0213",X"0198",X"0232",X"027C",X"034C",X"0400",X"04DA",X"05DA",X"06B9",X"06F0",X"0726",X"085A",X"0809",X"08EE",X"08F2",
		X"08B4",X"08A7",X"096D",X"0A8D",X"0B42",X"0B88",X"0D04",X"0DD8",X"0DB0",X"0E00",X"0ECF",X"0E1C",X"0D08",X"0CA3",X"0BB9",X"0A16",
		X"0857",X"07C2",X"071A",X"06C2",X"0610",X"0577",X"0588",X"05FC",X"05D7",X"054F",X"05C7",X"0572",X"0463",X"031D",X"02D6",X"025C",
		X"0180",X"00A0",X"004C",X"FFFB",X"FFAE",X"0042",X"002C",X"FF3A",X"0051",X"0112",X"FFCC",X"FE5A",X"FEA5",X"FF2D",X"FDDD",X"FCB8",
		X"FC89",X"FCC1",X"FB65",X"FBB4",X"FC82",X"FC11",X"FBA6",X"FC30",X"FBA4",X"FBBF",X"FCF9",X"FCF4",X"FC1D",X"FBF5",X"FC5D",X"FBF9",
		X"FC0B",X"FCD5",X"FD91",X"FCD8",X"FC8D",X"FDB7",X"FE0C",X"FEDD",X"FF32",X"FF33",X"FF4E",X"FEB6",X"FEEF",X"FF6E",X"FE57",X"FD95",
		X"FDA4",X"FD1A",X"FC32",X"FA88",X"FB2A",X"FB5B",X"FAA4",X"F9D1",X"FAB0",X"FA99",X"FA72",X"FAE4",X"FB1A",X"FBA3",X"FB16",X"FAEF",
		X"FAAD",X"FA6D",X"FA64",X"FA99",X"F9C1",X"F9F7",X"F99A",X"FA1E",X"F9B1",X"F9EF",X"FACB",X"FA97",X"FA6E",X"FAA0",X"FB87",X"F9BF",
		X"FB80",X"FAC7",X"FC48",X"FA22",X"FCBC",X"FBE4",X"FD49",X"FCC7",X"FEDF",X"FE56",X"FEFA",X"00A8",X"007A",X"01B8",X"015C",X"0389",
		X"01AC",X"0253",X"0307",X"0348",X"0264",X"03B1",X"022F",X"0444",X"01E5",X"0576",X"02F9",X"0608",X"0422",X"0644",X"0527",X"06D0",
		X"068D",X"0632",X"0764",X"04F8",X"0803",X"03A2",X"075D",X"04F3",X"0687",X"054A",X"04C0",X"05F3",X"055E",X"04D0",X"05E0",X"0456",
		X"04F0",X"04DB",X"0312",X"0513",X"029F",X"04BD",X"0356",X"01F1",X"048A",X"02D3",X"0289",X"042F",X"014A",X"03F4",X"01BC",X"022B",
		X"038E",X"010C",X"0288",X"0251",X"01A9",X"02CE",X"01FB",X"00FC",X"04B2",X"FF37",X"02E8",X"030D",X"FEE2",X"03EC",X"0169",X"FFB6",
		X"017D",X"00A2",X"FF43",X"FFF5",X"FF60",X"FE51",X"FEA6",X"FDF0",X"FC19",X"FDF4",X"FE93",X"FBBF",X"FE4C",X"FD69",X"FD79",X"FEAC",
		X"FCAF",X"FF51",X"FE7B",X"FCCC",X"FF87",X"FE0F",X"FC4A",X"FEDB",X"FED4",X"FCA7",X"FD98",X"FF90",X"FDB0",X"FC4E",X"0040",X"FF87",
		X"FC88",X"FF6C",X"0144",X"FC86",X"FE0B",X"01F9",X"FE0E",X"FCB0",X"FFF7",X"002B",X"FBC9",X"FE44",X"0075",X"FC23",X"FE16",X"0032",
		X"FCDD",X"FE2C",X"FED7",X"FDE3",X"FD70",X"FE0B",X"FF3F",X"FD21",X"FC6F",X"FEA0",X"FD84",X"FBCE",X"FDE8",X"FF83",X"FD00",X"FC8D",
		X"FEB3",X"FF68",X"FD29",X"FCCA",X"0057",X"FD8E",X"FB0A",X"FD3A",X"FF7D",X"FCB4",X"F9C5",X"FEB5",X"FFF1",X"FB17",X"FC16",X"0115",
		X"FF3E",X"FB61",X"FF9E",X"0231",X"FCE8",X"FCC1",X"025E",X"FFB8",X"FBAE",X"FFF6",X"02F9",X"FCB8",X"FC0B",X"038F",X"0111",X"FBFA",
		X"FFA6",X"0461",X"FF06",X"FD02",X"02DE",X"0361",X"FD68",X"FE8C",X"04FE",X"0021",X"FD08",X"019C",X"03D8",X"FE60",X"FF36",X"04B5",
		X"033F",X"FE89",X"01F7",X"064E",X"00D5",X"FF1E",X"03FC",X"058E",X"FF2C",X"FF52",X"0551",X"0494",X"FEE9",X"0100",X"069F",X"03EC",
		X"FF15",X"0250",X"057B",X"01B2",X"FE2D",X"0218",X"02DD",X"FDA4",X"FDA0",X"02A2",X"017A",X"FDF0",X"FFC5",X"02C6",X"02E1",X"0155",
		X"0388",X"0411",X"03C3",X"04D2",X"0631",X"03F2",X"046E",X"0642",X"05BB",X"03FE",X"050D",X"06E1",X"061E",X"059E",X"05AC",X"06D9",
		X"0656",X"07AC",X"05F6",X"04C8",X"064C",X"07A8",X"056C",X"02A1",X"04A8",X"0707",X"0498",X"0127",X"03E0",X"064B",X"03CF",X"015D",
		X"03C2",X"058F",X"02B4",X"0155",X"02C2",X"0215",X"00B4",X"001B",X"FFFB",X"FEAE",X"FE2F",X"FE43",X"FD55",X"FC37",X"FD3B",X"FD21",
		X"FABF",X"FA3B",X"FB34",X"FAB0",X"F854",X"F80C",X"F874",X"F772",X"F73A",X"F644",X"F68E",X"F6AB",X"F616",X"F505",X"F5E4",X"F5E9",
		X"F529",X"F57F",X"F568",X"F5CA",X"F66A",X"F5E5",X"F544",X"F6B7",X"F795",X"F73A",X"F4CF",X"F766",X"F93A",X"F761",X"F654",X"F8F8",
		X"F9FA",X"F8B2",X"F95C",X"FA13",X"FA0B",X"FA10",X"FB6B",X"FA6D",X"FA24",X"FB51",X"FC95",X"FBD7",X"FB38",X"FCE7",X"FEC3",X"FE66",
		X"FDC6",X"FED8",X"FFE7",X"0044",X"FED5",X"0018",X"0127",X"FF80",X"FFA4",X"0068",X"0093",X"00B6",X"0162",X"0164",X"015A",X"00E8",
		X"023D",X"043D",X"0266",X"031A",X"0479",X"05AB",X"04BC",X"04F2",X"0642",X"072C",X"06F7",X"06FB",X"076B",X"0805",X"0948",X"089B",
		X"0808",X"0844",X"0A25",X"08F0",X"07A3",X"086F",X"09F6",X"087C",X"079C",X"095C",X"0AA9",X"0936",X"09B5",X"0BBD",X"0AEF",X"0A91",
		X"0BB1",X"0C3F",X"0A9D",X"0AA4",X"0BBC",X"0ABA",X"08FF",X"09CD",X"09BF",X"08D4",X"07B0",X"0856",X"085B",X"071E",X"0688",X"06DD",
		X"077C",X"0697",X"053D",X"0531",X"0515",X"0417",X"0391",X"029E",X"01F1",X"00D5",X"0140",X"009D",X"FF5D",X"FF8D",X"00B7",X"FF80",
		X"FDF3",X"FEFF",X"FFFD",X"FEFC",X"FD4F",X"FDE3",X"FE56",X"FD3B",X"FC5B",X"FB62",X"FB64",X"FB74",X"FB14",X"FA5C",X"FA1E",X"FA66",
		X"FAD4",X"F952",X"F880",X"F8D9",X"F829",X"F6E8",X"F5C1",X"F5CE",X"F4F9",X"F42F",X"F498",X"F4D9",X"F469",X"F4A1",X"F61E",X"F614",
		X"F58E",X"F660",X"F714",X"F674",X"F57A",X"F65C",X"F6CD",X"F58F",X"F423",X"F5BF",X"F68B",X"F4DE",X"F560",X"F700",X"F730",X"F6F3",
		X"F795",X"F921",X"F93A",X"F9B7",X"F9F3",X"FA48",X"FA01",X"FA77",X"FA7B",X"FA3E",X"FA8E",X"FB42",X"FBF6",X"FB58",X"FCBE",X"FDB1",
		X"FE70",X"FE9E",X"FFD8",X"FFF8",X"0096",X"00E8",X"00F1",X"00DD",X"0148",X"0132",X"0099",X"0112",X"0180",X"01C3",X"0270",X"0348",
		X"03DA",X"043C",X"04ED",X"0534",X"060E",X"067F",X"0633",X"072F",X"0669",X"0717",X"070A",X"0748",X"0754",X"07CA",X"0859",X"0914",
		X"0A23",X"0A9B",X"0B0E",X"0C73",X"0D68",X"0CC4",X"0C9C",X"0C85",X"0C36",X"0B0B",X"0A74",X"0A01",X"091F",X"0758",X"074A",X"06F9",
		X"06F3",X"072E",X"0702",X"0656",X"061F",X"06B5",X"067E",X"055D",X"0492",X"0460",X"036E",X"01EE",X"00FD",X"0181",X"010B",X"FFB7",
		X"FF76",X"FFEA",X"007B",X"0128",X"009F",X"0083",X"00BA",X"00A6",X"FF56",X"FED9",X"FEC1",X"FE38",X"FD07",X"FC37",X"FC57",X"FC46",
		X"FC07",X"FC0E",X"FBDD",X"FBDF",X"FC46",X"FC0A",X"FC56",X"FCCF",X"FD16",X"FD1B",X"FCAF",X"FD1D",X"FD70",X"FD86",X"FDA3",X"FE1E",
		X"FE9A",X"FEA0",X"FF64",X"FF52",X"FFB2",X"0011",X"005F",X"00A4",X"FFC5",X"FF50",X"FF1D",X"FECF",X"FE4F",X"FE1C",X"FD35",X"FD0A",
		X"FC06",X"FBDA",X"FC59",X"FC6F",X"FC3A",X"FC23",X"FBFD",X"FC2E",X"FC17",X"FBF2",X"FC75",X"FBE1",X"FBFD",X"FB1E",X"FABE",X"FA8A",
		X"FAE8",X"FAEB",X"FA22",X"FA04",X"FA4B",X"FA7D",X"F9E0",X"FA0D",X"F9DB",X"FA7D",X"F944",X"FA99",X"F990",X"FA63",X"F93E",X"FAA5",
		X"F991",X"FAD5",X"FAC5",X"FC52",X"FC18",X"FC51",X"FE25",X"FDE1",X"0026",X"FF14",X"0163",X"0032",X"0153",X"008C",X"017C",X"0120",
		X"0144",X"FF76",X"016E",X"FF4B",X"01B1",X"FFEC",X"0206",X"007A",X"031D",X"0209",X"02F5",X"039B",X"0446",X"0508",X"0315",X"068F",
		X"031F",X"06CD",X"0334",X"0654",X"04C2",X"05AF",X"05EF",X"04C1",X"060E",X"0613",X"0523",X"05D0",X"0540",X"04AA",X"0591",X"0351",
		X"0543",X"030B",X"0375",X"0460",X"022B",X"047A",X"0475",X"030C",X"058D",X"02E5",X"04FC",X"04AB",X"0248",X"0473",X"02BD",X"0285",
		X"027E",X"0111",X"0220",X"0266",X"FF55",X"0440",X"0078",X"003B",X"045F",X"FFC4",X"0319",X"0330",X"009F",X"030A",X"022B",X"0000",
		X"00AF",X"010E",X"FEA1",X"FEA3",X"FFAA",X"FDFC",X"FD84",X"FEE2",X"FD59",X"FE9B",X"FF04",X"FDD0",X"FFA4",X"FE1B",X"FF2A",X"008B",
		X"FE17",X"FF2F",X"0024",X"FDB0",X"FF37",X"0034",X"FE83",X"FD8D",X"FFB3",X"0006",X"FCB9",X"FEC2",X"0147",X"FCFC",X"FCCC",X"00D8",
		X"FDC6",X"FB2E",X"FF94",X"FF01",X"FBDB",X"FD8F",X"003D",X"FD2F",X"FC13",X"00DB",X"FDD3",X"FCB1",X"0101",X"FF87",X"FF87",X"016F",
		X"0235",X"01A7",X"013D",X"039E",X"026C",X"FE70",X"FE62",X"FFC5",X"FC98",X"FB01",X"FB68",X"FA68",X"F878",X"F906",X"FB47",X"FB0E",
		X"F8EF",X"FB47",X"FCB6",X"FA0A",X"FA9B",X"FC9F",X"FD92",X"F90F",X"F9A5",X"FD0B",X"FAB0",X"F956",X"FCD1",X"FEDE",X"FB16",X"FBD2",
		X"0174",X"FFC4",X"FC54",X"01E7",X"02FA",X"FDB9",X"FD5F",X"033D",X"0173",X"FC99",X"0129",X"037F",X"FE69",X"FED0",X"04C0",X"03AF",
		X"FEC7",X"0266",X"0649",X"01FA",X"FF84",X"0646",X"06D0",X"01AF",X"03D3",X"07DD",X"0586",X"0298",X"06D2",X"0911",X"0605",X"04B2",
		X"08AF",X"07C7",X"05A5",X"065E",X"08EF",X"0759",X"047F",X"05FE",X"0677",X"04C2",X"0311",X"0519",X"0454",X"01C4",X"014F",X"0284",
		X"019E",X"000F",X"00D2",X"01B6",X"FFEC",X"FE93",X"0074",X"005E",X"FF25",X"FED2",X"FF97",X"FEBF",X"FD43",X"FEAC",X"FEAF",X"FD10",
		X"FD59",X"FEE6",X"FD27",X"FB21",X"FDB2",X"FE1D",X"FC90",X"FC5D",X"FDEB",X"FCF5",X"FBF9",X"FCB6",X"FE12",X"FC84",X"FBC1",X"FE5D",
		X"FDFD",X"FCC8",X"FDA0",X"FF24",X"FEE8",X"FDD2",X"FF70",X"0083",X"FF05",X"FEC1",X"0097",X"FFE0",X"FE68",X"FEEB",X"FF69",X"FDC1",
		X"FCC0",X"FE9A",X"FDE9",X"FD16",X"FDDC",X"FFA8",X"FE7D",X"FD1A",X"FEB9",X"FF2F",X"FDAF",X"FDF1",X"FEB3",X"FE1F",X"FDA8",X"FE4E",
		X"FF9B",X"FEE6",X"FF61",X"006D",X"FFD1",X"FF1E",X"FF56",X"FFAA",X"FFB8",X"FF3E",X"FF01",X"FFF9",X"FF67",X"FE29",X"FFD8",X"0138",
		X"0021",X"0046",X"0128",X"015F",X"0092",X"00DE",X"0209",X"0089",X"FFC7",X"0097",X"0025",X"FF07",X"003C",X"00F9",X"FFA4",X"002F",
		X"0183",X"0120",X"007A",X"01F5",X"0220",X"0179",X"0164",X"01C9",X"0209",X"0176",X"0126",X"010C",X"00C7",X"0051",X"FFD3",X"FF55",
		X"0011",X"FF9C",X"FF20",X"007B",X"004A",X"0034",X"00DE",X"014D",X"01BB",X"01A5",X"01CF",X"022B",X"01AF",X"0164",X"02B2",X"0143",
		X"014D",X"0210",X"01A2",X"011C",X"0134",X"0233",X"0178",X"0120",X"014C",X"0197",X"0100",X"00DC",X"0126",X"00E1",X"005E",X"0088",
		X"0058",X"FF7C",X"FEF5",X"FFE6",X"FFED",X"FE72",X"FF13",X"0016",X"FF7F",X"FE4F",X"FFBF",X"FFE9",X"FEB0",X"FE87",X"FEE5",X"FE7F",
		X"FD59",X"FE18",X"FDC9",X"FCCE",X"FD1F",X"FDBD",X"FDD9",X"FD4D",X"FE0C",X"FEED",X"FE59",X"FE53",X"FEB6",X"FEF9",X"FE0F",X"FDC1",
		X"FE1E",X"FE2F",X"FD9B",X"FDBD",X"FE72",X"FEE3",X"FE7E",X"FF21",X"0072",X"00DF",X"00A1",X"00E1",X"0185",X"0147",X"012C",X"01BC",
		X"01AB",X"011B",X"0130",X"0164",X"015B",X"016B",X"01BE",X"01A9",X"0173",X"015E",X"01D8",X"0198",X"0191",X"0217",X"0257",X"0218",
		X"0213",X"0288",X"01D6",X"0212",X"02BD",X"023B",X"0203",X"01EC",X"026D",X"0259",X"01D0",X"0280",X"02F7",X"02AA",X"01FD",X"0239",
		X"02EF",X"02BB",X"01DA",X"0184",X"0247",X"0130",X"00E7",X"01CB",X"00F4",X"00DA",X"0163",X"0139",X"0131",X"016A",X"01A4",X"01B2",
		X"0102",X"0148",X"0181",X"006E",X"FFED",X"FFFC",X"FFDE",X"FF66",X"FF12",X"FF73",X"FEE8",X"FE93",X"FF1E",X"FE96",X"FE24",X"FE77",
		X"FE8C",X"FDBF",X"FE35",X"FE66",X"FDAE",X"FD70",X"FD87",X"FD48",X"FCAA",X"FC89",X"FC58",X"FBD3",X"FBB1",X"FBA5",X"FB68",X"FB98",
		X"FC02",X"FBF9",X"FC17",X"FBF6",X"FC6B",X"FC9D",X"FCE7",X"FD3E",X"FCD5",X"FCDE",X"FCA3",X"FD06",X"FCC9",X"FCF1",X"FD1D",X"FD43",
		X"FD2D",X"FD7C",X"FDF3",X"FDC8",X"FD8E",X"FDB8",X"FD3D",X"FD6E",X"FD38",X"FCC7",X"FD3C",X"FD6D",X"FDAE",X"FD45",X"FD8D",X"FE17",
		X"FE9A",X"FE4C",X"FF3E",X"FFD9",X"FF5C",X"FF9A",X"FFF8",X"0026",X"0054",X"0099",X"0103",X"008A",X"003E",X"0127",X"00B8",X"008E",
		X"00F0",X"0135",X"00F0",X"0184",X"0212",X"01E0",X"020A",X"01F1",X"0227",X"0250",X"020D",X"01CF",X"01CB",X"01BD",X"0237",X"0269",
		X"0252",X"030B",X"0395",X"036B",X"0413",X"046F",X"0489",X"04B0",X"046D",X"0433",X"04C2",X"0478",X"045A",X"0493",X"04A7",X"04F9",
		X"04B4",X"0528",X"051B",X"04DD",X"04B5",X"04D1",X"043A",X"0408",X"03D2",X"0319",X"0347",X"0262",X"02AA",X"0327",X"0300",X"036E",
		X"039D",X"037E",X"037D",X"037F",X"0324",X"02D0",X"0259",X"01C4",X"018E",X"0167",X"012D",X"011C",X"00AA",X"004D",X"0090",X"0046",
		X"0062",X"FFF9",X"FFB0",X"FF7C",X"FEBC",X"FE9D",X"FE7D",X"FE15",X"FE48",X"FE4E",X"FDD4",X"FE95",X"FEA4",X"FE7A",X"FE93",X"FE2D",
		X"FEB7",X"FDF8",X"FDB5",X"FDC6",X"FD66",X"FD6D",X"FCEC",X"FCC8",X"FC37",X"FC39",X"FB9C",X"FB70",X"FB6E",X"FB90",X"FB46",X"FB45",
		X"FBC9",X"FB64",X"FC1C",X"FBF7",X"FB98",X"FBD5",X"FBCF",X"FBB1",X"FB56",X"FB63",X"FB4B",X"FB24",X"FB42",X"FBC3",X"FB9E",X"FB86",
		X"FBF8",X"FC31",X"FC5E",X"FCA7",X"FC69",X"FCA9",X"FCF9",X"FD02",X"FD7F",X"FD94",X"FDA1",X"FE20",X"FE9C",X"FF28",X"FF40",X"FF68",
		X"FFCE",X"FFC9",X"FFD4",X"0022",X"0068",X"FFEE",X"FFC0",X"005B",X"0040",X"FFFF",X"002F",X"00B3",X"00E8",X"00E3",X"00C8",X"0145",
		X"0171",X"016C",X"01A9",X"0194",X"01BC",X"01BA",X"01C9",X"01E2",X"01E3",X"0233",X"0252",X"0201",X"022B",X"028B",X"0258",X"024B",
		X"0256",X"02CC",X"029C",X"026F",X"02DE",X"026F",X"02BD",X"0300",X"02D9",X"0332",X"035D",X"02E6",X"0333",X"030F",X"0365",X"0377",
		X"02FE",X"0399",X"03DC",X"0384",X"0395",X"041C",X"0435",X"03B3",X"0428",X"0506",X"04FF",X"046C",X"04AB",X"04A1",X"03CF",X"0373",
		X"0367",X"02F4",X"0255",X"021E",X"0233",X"01D7",X"01C9",X"0220",X"0226",X"0206",X"024E",X"027A",X"0231",X"01DE",X"01B3",X"0148",
		X"009F",X"0085",X"0039",X"0025",X"FFBF",X"FFDC",X"FFC0",X"FFCF",X"FFC5",X"0019",X"0061",X"004D",X"0001",X"0040",X"FFED",X"FF97",
		X"FFA6",X"FEFC",X"FE67",X"FDAC",X"FDD9",X"FE02",X"FDE3",X"FD53",X"FD97",X"FE07",X"FDD8",X"FD8C",X"FDA1",X"FD5B",X"FD3F",X"FD04",
		X"FCAE",X"FC45",X"FB94",X"FB8A",X"FAD2",X"FAFC",X"FB16",X"FB06",X"FB0C",X"FB5C",X"FBF7",X"FC28",X"FC08",X"FC33",X"FC45",X"FC01",
		X"FBCC",X"FB70",X"FB54",X"FAD9",X"FAD1",X"FA8B",X"FA70",X"FAFC",X"FAD7",X"FAF8",X"FBAD",X"FC2F",X"FBFC",X"FBE4",X"FBF8",X"FC21",
		X"FBD0",X"FB94",X"FB86",X"FB13",X"FB0F",X"FAC1",X"FB00",X"FB46",X"FBB4",X"FB94",X"FBBA",X"FC79",X"FD04",X"FD35",X"FD64",X"FDBF",
		X"FE09",X"FE9E",X"FE4E",X"FE5B",X"FF1C",X"FED9",X"FE8F",X"FEF1",X"FF83",X"FF99",X"FFB9",X"0009",X"00B9",X"00FB",X"0147",X"017C",
		X"017C",X"0229",X"024C",X"0275",X"029E",X"02C4",X"0326",X"0375",X"0381",X"041B",X"048D",X"0487",X"050E",X"055F",X"0593",X"057C",
		X"061F",X"0674",X"0611",X"06B0",X"06CB",X"0717",X"06E3",X"06F5",X"0729",X"074F",X"0759",X"072A",X"0724",X"0730",X"0790",X"06E9",
		X"06C6",X"06DD",X"0703",X"06C1",X"0693",X"072B",X"0701",X"0659",X"06A5",X"06D3",X"06D3",X"0691",X"0603",X"064E",X"0670",X"063E",
		X"05AD",X"05A0",X"0562",X"04D6",X"0404",X"0444",X"0418",X"02AA",X"0273",X"0252",X"019E",X"00E5",X"00AF",X"0015",X"FF51",X"FF19",
		X"FF07",X"FE9A",X"FE12",X"FDEA",X"FD95",X"FD2D",X"FCE8",X"FCD2",X"FBF1",X"FB68",X"FB8B",X"FAE5",X"FA60",X"FA58",X"FA4B",X"F9E4",
		X"F9CA",X"F9E6",X"F9E4",X"F9EB",X"F9B1",X"F991",X"F9A7",X"F9B7",X"F986",X"F8E6",X"F8C1",X"F908",X"F8FF",X"F8AA",X"F849",X"F882",
		X"F8ED",X"F8B4",X"F882",X"F8D8",X"F8C3",X"F8FF",X"F905",X"F928",X"F993",X"F9B8",X"F992",X"F9DD",X"FA3A",X"FA4C",X"FA6F",X"FA88",
		X"FB08",X"FB60",X"FBC5",X"FC2C",X"FCE2",X"FCF0",X"FCEF",X"FD48",X"FDA2",X"FD9A",X"FD61",X"FD72",X"FD7B",X"FDB1",X"FE08",X"FDCA",
		X"FE30",X"FF0B",X"FF1A",X"FF3C",X"FFDE",X"00A8",X"0099",X"00CD",X"01A5",X"01D2",X"01DC",X"0254",X"02CF",X"0318",X"03D9",X"0453",
		X"048F",X"0556",X"0640",X"0694",X"06D7",X"077E",X"07D4",X"07E7",X"07F0",X"0861",X"0865",X"0842",X"0831",X"0863",X"0870",X"084E",
		X"0848",X"07D3",X"0807",X"0839",X"07E0",X"0773",X"0749",X"0777",X"070F",X"064D",X"065C",X"063A",X"0593",X"055A",X"054A",X"051A",
		X"0521",X"04D1",X"046A",X"0474",X"0427",X"03F7",X"03C0",X"0338",X"02FD",X"0262",X"01E2",X"0182",X"0106",X"00B8",X"0073",X"FFE1",
		X"FFDF",X"FFD2",X"FF9F",X"FF8E",X"FF5A",X"FFA6",X"FF9E",X"FEEA",X"FE81",X"FE62",X"FE29",X"FD90",X"FCFD",X"FCD1",X"FCE1",X"FC6A",
		X"FBB4",X"FBEF",X"FC32",X"FBAD",X"FB7D",X"FB97",X"FB71",X"FB44",X"FB1B",X"FB3A",X"FAE1",X"FAE6",X"FAE6",X"FA9F",X"FAAA",X"FACB",
		X"FB2B",X"FB0A",X"FAF6",X"FB6F",X"FB79",X"FB74",X"FB5D",X"FBAD",X"FB32",X"FB1B",X"FB0E",X"FADE",X"FAEB",X"FB3C",X"FB2F",X"FB54",
		X"FBB2",X"FB80",X"FB9B",X"FBB3",X"FBEA",X"FBD1",X"FC53",X"FC60",X"FC1D",X"FC83",X"FCC8",X"FD00",X"FD3A",X"FD6B",X"FDA1",X"FDBC",
		X"FE0C",X"FE27",X"FE82",X"FEA8",X"FEB9",X"FF10",X"FFAF",X"FFEA",X"FFD3",X"FFDA",X"000D",X"FFD6",X"FFE4",X"007F",X"0045",X"0017",
		X"0087",X"00CF",X"00F8",X"0101",X"0118",X"01A2",X"01C1",X"01CC",X"0221",X"0262",X"0244",X"0270",X"02E5",X"031F",X"0336",X"034A",
		X"032E",X"032B",X"0362",X"0327",X"02DD",X"02D3",X"02B3",X"0270",X"0255",X"028B",X"02C1",X"02A7",X"0285",X"02C2",X"02B2",X"029E",
		X"026F",X"025D",X"0224",X"01E5",X"018B",X"0159",X"0161",X"017C",X"0166",X"0189",X"01B7",X"0203",X"025E",X"01F4",X"020A",X"0225",
		X"01DD",X"01AF",X"019D",X"0195",X"0154",X"0113",X"0166",X"019C",X"0165",X"016D",X"01E8",X"01CA",X"0180",X"01CF",X"01AF",X"0131",
		X"00CC",X"00E4",X"00EC",X"007C",X"005A",X"005B",X"0065",X"003B",X"0058",X"0070",X"0029",X"FFCB",X"FFCC",X"FFF4",X"FFE0",X"FFD2",
		X"0015",X"FFFA",X"FFD7",X"002D",X"006E",X"0040",X"004F",X"005F",X"003A",X"0070",X"0065",X"007C",X"0084",X"00A7",X"00BA",X"00D2",
		X"00F6",X"00B1",X"0056",X"0068",X"0042",X"FFF7",X"FFCE",X"FF81",X"FF15",X"FED2",X"FF23",X"FF33",X"FE98",X"FEC0",X"FEF2",X"FE99",
		X"FEA7",X"FEDA",X"FEF7",X"FE7F",X"FEA1",X"FED8",X"FEB2",X"FE4E",X"FE2D",X"FDEA",X"FD6C",X"FD69",X"FD60",X"FD49",X"FD1F",X"FD97",
		X"FDCB",X"FDA6",X"FDDD",X"FE39",X"FE48",X"FE57",X"FEDA",X"FEFB",X"FEE6",X"FF04",X"FF11",X"FED5",X"FEDD",X"FF18",X"FF1B",X"FF05",
		X"FEF9",X"FEC8",X"FE95",X"FEE9",X"FEE3",X"FE75",X"FEBF",X"FEC8",X"FE8C",X"FE95",X"FE91",X"FE92",X"FE52",X"FE38",X"FEBC",X"FEE6",
		X"FEEE",X"FF2E",X"FF71",X"FF8C",X"FFBA",X"FFF4",X"FFC8",X"FFF4",X"FFF9",X"0028",X"0067",X"008D",X"00D1",X"00F0",X"010F",X"0124",
		X"013D",X"014C",X"0127",X"00E9",X"00C5",X"009C",X"0075",X"0050",X"003D",X"0071",X"001F",X"0018",X"0082",X"0095",X"0090",X"00E2",
		X"0125",X"017A",X"01E0",X"022E",X"028B",X"02B2",X"02EF",X"0329",X"0325",X"032D",X"0349",X"0315",X"02FA",X"02E9",X"02C2",X"0295",
		X"0286",X"0274",X"025A",X"0248",X"023E",X"0250",X"0287",X"02AB",X"02A3",X"027B",X"026B",X"028A",X"025B",X"01F9",X"01BF",X"01B7",
		X"0170",X"0152",X"013E",X"010B",X"00F5",X"00CA",X"00A2",X"007A",X"0065",X"0018",X"FF7E",X"FF89",X"FFC5",X"FFA0",X"FF72",X"FF85",
		X"FF90",X"FF7F",X"FF80",X"FF9F",X"FF98",X"FF86",X"FFA3",X"FF5F",X"FF22",X"FF33",X"FF29",X"FEE2",X"FEB2",X"FEC3",X"FEA6",X"FE64",
		X"FE6A",X"FE5D",X"FE43",X"FE25",X"FE16",X"FDD7",X"FE13",X"FDFB",X"FE09",X"FDFF",X"FDE9",X"FDF3",X"FDB5",X"FD75",X"FD6E",X"FD9B",
		X"FD57",X"FD2F",X"FD79",X"FD9B",X"FDC8",X"FDE6",X"FDF1",X"FE2A",X"FE21",X"FE05",X"FDA8",X"FD9A",X"FD81",X"FD67",X"FD3E",X"FD30",
		X"FD8D",X"FDB0",X"FDE7",X"FE2D",X"FE99",X"FEEC",X"FED7",X"FF23",X"FF1F",X"FEDD",X"FEDC",X"FF0E",X"FF15",X"FEF9",X"FF03",X"FF34",
		X"FF2D",X"FF11",X"FF59",X"FF23",X"FEEE",X"FF30",X"FF3E",X"FF5B",X"FFA3",X"FF93",X"FFA8",X"FFED",X"002B",X"0054",X"00AD",X"00E2",
		X"010C",X"0124",X"0135",X"0162",X"018D",X"01AE",X"017C",X"0170",X"0182",X"0184",X"014F",X"0161",X"0183",X"015D",X"014C",X"0180",
		X"0193",X"014F",X"0123",X"011E",X"013A",X"0146",X"0156",X"017D",X"0155",X"0181",X"01B0",X"0199",X"016E",X"01A7",X"01AA",X"0112",
		X"00DB",X"011D",X"00C6",X"0064",X"00AD",X"00D3",X"00A6",X"0099",X"00F6",X"013B",X"00E8",X"0128",X"016D",X"0122",X"0101",X"0108",
		X"00AE",X"001E",X"003F",X"006A",X"0035",X"FFC6",X"FFE6",X"0044",X"003C",X"0012",X"0042",X"0056",X"0039",X"006B",X"0053",X"0055",
		X"0016",X"0014",X"0030",X"002B",X"002B",X"0013",X"0027",X"FFC5",X"FFC9",X"000E",X"FFF4",X"FF87",X"FF8E",X"FFAB",X"FFD8",X"FFB5",
		X"FFB7",X"FFB7",X"FFC3",X"FFD3",X"FFFC",X"0038",X"0023",X"0079",X"00CA",X"00EB",X"011A",X"0133",X"012E",X"0120",X"011D",X"014D",
		X"0120",X"00FA",X"00CD",X"0095",X"004B",X"004F",X"0016",X"0003",X"0020",X"0014",X"000F",X"0038",X"0068",X"0079",X"005F",X"0039",
		X"004D",X"0034",X"0020",X"FFF0",X"FFCF",X"FF99",X"FF5F",X"FF81",X"FF84",X"FF74",X"FF48",X"FF3F",X"FF98",X"FF75",X"FF83",X"FF78",
		X"FF56",X"FF20",X"FF08",X"FEFD",X"FECB",X"FE7C",X"FE5A",X"FE59",X"FE6E",X"FE79",X"FE7A",X"FE9B",X"FE9C",X"FE84",X"FEBB",X"FEFE",
		X"FEC9",X"FE7B",X"FE76",X"FE78",X"FE43",X"FE38",X"FE33",X"FE48",X"FE12",X"FE3E",X"FEB4",X"FF00",X"FEE7",X"FEF1",X"FEFF",X"FEF6",
		X"FF08",X"FEEF",X"FED8",X"FECA",X"FEA6",X"FEAF",X"FEF2",X"FF26",X"FF17",X"FF13",X"FF34",X"FF64",X"FFB0",X"0001",X"0009",X"0008",
		X"0031",X"0025",X"0007",X"FFE7",X"001A",X"0029",X"000C",X"003E",X"0055",X"0064",X"007D",X"00BD",X"00F7",X"0165",X"018F",X"0186",
		X"01CB",X"024E",X"026B",X"0231",X"026C",X"02A1",X"027A",X"02B1",X"02E3",X"02C2",X"028F",X"027A",X"0276",X"0291",X"02CF",X"02FF",
		X"02CA",X"0298",X"02CC",X"02C2",X"029C",X"0294",X"0290",X"024F",X"0272",X"0252",X"0231",X"023E",X"0212",X"01DE",X"01CB",X"01F5",
		X"01EC",X"018F",X"0173",X"017F",X"0148",X"00D5",X"00BE",X"0090",X"0058",X"0043",X"000F",X"FFE4",X"FFDB",X"0002",X"FFDE",X"FFD3",
		X"0002",X"FFDF",X"FF90",X"FF6D",X"FF7F",X"FF55",X"FEF6",X"FED1",X"FE6D",X"FE29",X"FDF4",X"FDD0",X"FDA6",X"FDBF",X"FDA9",X"FD9F",
		X"FDBC",X"FDFC",X"FE09",X"FDDC",X"FDFD",X"FE05",X"FDE3",X"FDB4",X"FE12",X"FE23",X"FDDA",X"FDD8",X"FE1C",X"FDE7",X"FDE1",X"FE3A",
		X"FE8D",X"FE9B",X"FE89",X"FEAE",X"FE8C",X"FEB5",X"FED2",X"FEC6",X"FEA0",X"FE9D",X"FE7F",X"FE36",X"FE03",X"FE0B",X"FDE7",X"FDC4",
		X"FD9B",X"FD99",X"FDA1",X"FD93",X"FDB4",X"FDCA",X"FE1D",X"FE3F",X"FE80",X"FE71",X"FE6E",X"FEB1",X"FF0E",X"FF05",X"FEF5",X"FF38",
		X"FF69",X"FF68",X"FF8A",X"0008",X"004C",X"004D",X"0050",X"009C",X"00C6",X"00B3",X"00B5",X"00DE",X"00F5",X"0103",X"010A",X"011D",
		X"0157",X"01A8",X"01E6",X"01D9",X"01CD",X"0201",X"020F",X"01F8",X"0246",X"0263",X"0222",X"01E5",X"021D",X"0248",X"0220",X"01EF",
		X"01D5",X"019A",X"019D",X"01AA",X"01A3",X"0186",X"0159",X"0179",X"018C",X"01A8",X"019E",X"01A3",X"017D",X"015B",X"0123",X"0118",
		X"00FC",X"0106",X"00FE",X"00D7",X"00BE",X"00AF",X"00C6",X"00CE",X"00BC",X"00C8",X"0098",X"0045",X"004D",X"001B",X"FFAD",X"FF62",
		X"FF63",X"FF1E",X"FEC6",X"FEAB",X"FE9D",X"FE41",X"FE05",X"FE03",X"FE11",X"FDEA",X"FE0D",X"FE2E",X"FE45",X"FE6D",X"FEB3",X"FEFE",
		X"FF49",X"FFA5",X"FFA8",X"FFB7",X"FFDA",X"FFE5",X"FFB9",X"FF94",X"FF99",X"FF85",X"FF5E",X"FF47",X"FF24",X"FF1F",X"FF52",X"FF5C",
		X"FF50",X"FF3B",X"FF45",X"FF76",X"FF2B",X"FF34",X"FF66",X"FF4A",X"FF48",X"FF61",X"FF88",X"FFEC",X"002B",X"0059",X"0057",X"0043",
		X"0059",X"008B",X"0073",X"0076",X"0064",X"0074",X"0067",X"007B",X"0087",X"0090",X"00C1",X"012C",X"014F",X"0173",X"019C",X"016D",
		X"0151",X"013A",X"0130",X"00EF",X"00EE",X"00D8",X"00A3",X"0082",X"0072",X"0054",X"000C",X"FFEA",X"FFDE",X"FF97",X"FF94",X"FFA6",
		X"FFCE",X"FFE8",X"FFCD",X"FFC0",X"FFD8",X"FFF3",X"0005",X"002B",X"0027",X"0001",X"0033",X"0035",X"0028",X"0037",X"007F",X"0092",
		X"003B",X"003C",X"0055",X"001B",X"0006",X"0014",X"FFF4",X"FFFA",X"0013",X"0030",X"004D",X"0089",X"00D1",X"00C3",X"00D4",X"0110",
		X"015B",X"0134",X"00F1",X"00C1",X"00BC",X"0096",X"003A",X"0018",X"FFFE",X"FFDF",X"FFBB",X"FFB1",X"FFC8",X"FFBD",X"FFBB",X"FFD7",
		X"FFDD",X"FFBF",X"FFB0",X"FFAE",X"FF97",X"FF79",X"FF89",X"FFB7",X"FFB7",X"FFCD",X"FFCA",X"FFD1",X"FFD6",X"FFC6",X"FFCE",X"FFB4",
		X"FF9B",X"FFC4",X"FFE9",X"FFC7",X"FF8A",X"FF92",X"FFCC",X"FF94",X"FF64",X"FF7E",X"FF70",X"FF60",X"FF7F",X"FF8B",X"FFB0",X"FFB5",
		X"FFD8",X"FFEA",X"FFFA",X"002F",X"001A",X"FFE6",X"FF82",X"FF52",X"FF48",X"FF3C",X"FF13",X"FEFF",X"FF26",X"FF54",X"FF8D",X"FFC8",
		X"FFE4",X"0019",X"0050",X"006E",X"0069",X"0083",X"0084",X"0040",X"FFF9",X"FFEC",X"FFE8",X"FFA6",X"FF79",X"FF5A",X"FF84",X"FF85",
		X"FF90",X"FFAA",X"FFC9",X"FFFB",X"003D",X"0081",X"0085",X"008C",X"0084",X"0089",X"007A",X"005E",X"0036",X"0029",X"0021",X"0023",
		X"001A",X"0048",X"007B",X"0094",X"00A7",X"00C4",X"00B8",X"0093",X"0081",X"008C",X"0071",X"0016",X"FFE7",X"FFDC",X"FFB5",X"FFCB",
		X"0000",X"0038",X"0076",X"00D9",X"011A",X"0147",X"015F",X"015A",X"014E",X"00FE",X"00BD",X"0068",X"FFF4",X"FFC8",X"FFB0",X"FFB8",
		X"FFB8",X"FFDE",X"FFED",X"0009",X"000C",X"0004",X"0025",X"FFEB",X"FFCB",X"FF93",X"FF95",X"FF9A",X"FFC8",X"FFA7",X"FF9B",X"FF75",
		X"FFA4",X"FFDD",X"FFCB",X"FFA3",X"FFCB",X"0003",X"0012",X"005E",X"0057",X"FFFA",X"FFAF",X"FFBF",X"FFA6",X"FF45",X"FF03",X"FF05",
		X"FEEF",X"FEF5",X"FF1D",X"FF69",X"FF61",X"FF68",X"FFB1",X"FFD1",X"FF9E",X"FF79",X"FF74",X"FF44",X"FF10",X"FEE4",X"FEA5",X"FE6F",
		X"FE82",X"FEC9",X"FED1",X"FEFA",X"FF26",X"FF65",X"FF70",X"FF85",X"FF69",X"FF74",X"FF98",X"FF5E",X"FF4F",X"FF3D",X"FF30",X"FF03",
		X"FF02",X"FF29",X"FF5C",X"FF50",X"FF60",X"FF44",X"FF93",X"FFCC",X"FFB2",X"FFA2",X"FFB0",X"FFAB",X"FF96",X"FFCE",X"FFDB",X"FFFC",
		X"000C",X"0006",X"FFE3",X"FFC2",X"FFA7",X"FF7E",X"FF1A",X"FF2F",X"FF60",X"FF17",X"FF17",X"FF49",X"FF90",X"FFB8",X"FFF0",X"0057",
		X"006B",X"005D",X"0088",X"0084",X"0058",X"0041",X"004F",X"002D",X"001D",X"003C",X"004B",X"FFF9",X"FFBE",X"FFFA",X"0011",X"0013",
		X"001E",X"0028",X"0075",X"009F",X"00D6",X"0121",X"016B",X"017C",X"0196",X"01C0",X"01CE",X"01B0",X"0188",X"016A",X"0158",X"017B",
		X"017E",X"0162",X"0156",X"0165",X"01A1",X"01D4",X"01D2",X"020A",X"0233",X"0242",X"0236",X"0239",X"0241",X"021E",X"0238",X"0260",
		X"0250",X"024A",X"0232",X"0205",X"01E4",X"01D2",X"0168",X"010A",X"00F9",X"00DE",X"008C",X"0045",X"002F",X"0045",X"0040",X"0042",
		X"0056",X"0023",X"0019",X"0014",X"000D",X"0010",X"FFE2",X"FFC7",X"FFF9",X"000E",X"0022",X"FFFF",X"FFCA",X"FFB7",X"FFB4",X"FF92",
		X"FF6C",X"FF59",X"FF7A",X"FF66",X"FF23",X"FF1C",X"FF21",X"FF1E",X"FEEA",X"FEC6",X"FEC5",X"FEB3",X"FE9F",X"FE90",X"FE8E",X"FE73",
		X"FE69",X"FE77",X"FE8A",X"FE84",X"FE75",X"FEA9",X"FE8D",X"FE8B",X"FE93",X"FE83",X"FE9E",X"FE9D",X"FEC0",X"FED5",X"FF07",X"FF08",
		X"FEBE",X"FE83",X"FE93",X"FE64",X"FE13",X"FE2D",X"FE61",X"FE9B",X"FEA2",X"FE9E",X"FEA4",X"FEF5",X"FF45",X"FF54",X"FF25",X"FF2F",
		X"FF1F",X"FF16",X"FF17",X"FEEE",X"FEDE",X"FE94",X"FE72",X"FE8B",X"FEB5",X"FEE4",X"FF0E",X"FF4E",X"FFA7",X"002A",X"0055",X"008F",
		X"00CE",X"0117",X"0175",X"016C",X"0173",X"017D",X"0166",X"013F",X"0136",X"013C",X"013F",X"013D",X"0166",X"019B",X"0196",X"01C2",
		X"01CB",X"01EB",X"01FD",X"0211",X"0204",X"0201",X"022A",X"01FD",X"01F5",X"01E4",X"01E2",X"01F2",X"0217",X"01DF",X"01B5",X"01A3",
		X"0190",X"017E",X"0145",X"011E",X"00E7",X"00DF",X"00DC",X"00DD",X"00DD",X"00D0",X"00C9",X"00EA",X"011A",X"0152",X"0152",X"0116",
		X"0104",X"00F9",X"00CA",X"00B7",X"0096",X"005B",X"003D",X"0020",X"0017",X"0016",X"0005",X"FFE6",X"FFE9",X"003A",X"0049",X"002E",
		X"000A",X"FFFE",X"0034",X"0070",X"0068",X"0072",X"0035",X"0005",X"FFCD",X"FFEC",X"FFF7",X"FFB7",X"FF8C",X"FF1B",X"FF36",X"FF49",
		X"FF42",X"FF2B",X"FF1B",X"FEF1",X"FEED",X"FEF2",X"FEE2",X"FEF3",X"FEFA",X"FEFC",X"FEE4",X"FEB0",X"FECC",X"FE9D",X"FE5D",X"FE50",
		X"FE19",X"FDF0",X"FD8C",X"FD55",X"FD5B",X"FD4F",X"FD56",X"FD84",X"FD89",X"FDAE",X"FDFF",X"FE0E",X"FE22",X"FE19",X"FE2A",X"FE2F",
		X"FE10",X"FE41",X"FE47",X"FE49",X"FE2D",X"FE1C",X"FE6B",X"FE7E",X"FE7E",X"FE96",X"FEA4",X"FEA7",X"FEB8",X"FEC5",X"FEE8",X"FEE7",
		X"FEE9",X"FEB5",X"FE96",X"FEAF",X"FEBB",X"FF0F",X"FF34",X"FF5D",X"FF76",X"FF83",X"FFCF",X"0004",X"0045",X"005E",X"007A",X"00C3",
		X"00D8",X"00DA",X"010F",X"0139",X"0122",X"0120",X"0151",X"0168",X"0156",X"0143",X"016C",X"0153",X"00E8",X"00D4",X"00BC",X"009C",
		X"009E",X"0084",X"006B",X"0077",X"007D",X"00C2",X"00EB",X"0101",X"0149",X"015F",X"0161",X"017A",X"0176",X"0179",X"0147",X"0118",
		X"0121",X"00E2",X"00EE",X"013E",X"0169",X"0148",X"0128",X"012F",X"013D",X"0122",X"011E",X"012B",X"0117",X"00F9",X"00F0",X"00CC",
		X"0079",X"0091",X"00E5",X"00BD",X"00A5",X"00E1",X"0108",X"00D9",X"00C4",X"00EA",X"0107",X"00FF",X"00F0",X"00E5",X"00D1",X"00E4",
		X"00F5",X"00FB",X"0134",X"0154",X"017A",X"0197",X"01A8",X"01EC",X"01EA",X"01D9",X"01BB",X"017D",X"013D",X"0118",X"00F2",X"00CB",
		X"00C5",X"00AD",X"00B0",X"0090",X"0076",X"0066",X"0035",X"0018",X"0000",X"FFCB",X"FF8C",X"FF39",X"FF22",X"FEE9",X"FE83",X"FE50",
		X"FE31",X"FE33",X"FE10",X"FDD5",X"FD96",X"FD9B",X"FD8C",X"FDB5",X"FD96",X"FD8E",X"FD7C",X"FD66",X"FD9D",X"FDBA",X"FD9F",X"FD52",
		X"FD3D",X"FD46",X"FD7C",X"FD9E",X"FDCC",X"FDB7",X"FDED",X"FE21",X"FE3D",X"FE71",X"FE7C",X"FE93",X"FE85",X"FE85",X"FEAA",X"FEAA",
		X"FE94",X"FE8A",X"FEC0",X"FED3",X"FF07",X"FF73",X"FFB9",X"FFAF",X"FFCC",X"FFDB",X"FFE0",X"FFAF",X"FF8A",X"FFB8",X"FFC0",X"FFE0",
		X"FFE2",X"FFF8",X"0009",X"0048",X"0098",X"00B9",X"00DE",X"0117",X"013E",X"0129",X"0152",X"0181",X"0176",X"015A",X"015E",X"017A",
		X"0142",X"0138",X"014A",X"015B",X"0148",X"015D",X"0150",X"0159",X"0169",X"0166",X"018C",X"0196",X"01A6",X"01A4",X"01A1",X"01B1",
		X"01F2",X"022A",X"0245",X"0237",X"025B",X"0293",X"0280",X"026E",X"0294",X"0277",X"024D",X"022F",X"0210",X"021C",X"020C",X"01ED",
		X"01E0",X"01B9",X"01BB",X"01B2",X"01B1",X"019B",X"019B",X"01AE",X"0190",X"0174",X"014F",X"0149",X"0123",X"010F",X"00E7",X"0099",
		X"006C",X"0058",X"003F",X"0026",X"0021",X"FFED",X"FFBE",X"FFBC",X"FF96",X"FF64",X"FF52",X"FF52",X"FF15",X"FEEC",X"FEE8",X"FED1",
		X"FECE",X"FEB3",X"FE96",X"FE4C",X"FE42",X"FE1A",X"FDE5",X"FDA9",X"FD65",X"FD5C",X"FD3B",X"FD12",X"FD18",X"FD26",X"FD56",X"FD6D",
		X"FD8E",X"FDF3",X"FE51",X"FE7C",X"FE81",X"FE6E",X"FE3F",X"FE1D",X"FDEA",X"FDE9",X"FDDB",X"FDDC",X"FDCB",X"FDED",X"FE3C",X"FEA6",
		X"FEBF",X"FECC",X"FEB8",X"FED4",X"FEDA",X"FEE1",X"FEE0",X"FEC5",X"FEBF",X"FEFA",X"FF42",X"FF51",X"FF87",X"FF98",X"FFD3",X"FFED",
		X"0023",X"003D",X"0037",X"003B",X"0050",X"0062",X"0041",X"004A",X"0052",X"0048",X"0051",X"0059",X"0044",X"0038",X"004E",X"004A",
		X"0048",X"0049",X"001B",X"0007",X"0023",X"004A",X"006C",X"0059",X"0065",X"0083",X"008A",X"009D",X"00BD",X"00E0",X"00FE",X"011C",
		X"0134",X"0141",X"0173",X"0183",X"0159",X"018A",X"0186",X"0165",X"014C",X"0108",X"00C0",X"00A3",X"00AA",X"0092",X"0079",X"0096",
		X"00CA",X"00B1",X"00DF",X"011D",X"0115",X"0108",X"010A",X"0131",X"0116",X"00F1",X"00AE",X"0062",X"0030",X"FFFD",X"FFA6",X"FF87",
		X"FF93",X"FF97",X"FFAC",X"FFB6",X"FFD6",X"FFE4",X"FFD6",X"FFDB",X"FFE9",X"FFDC",X"FF85",X"FF2B",X"FEFE",X"FEE5",X"FEC0",X"FE9D",
		X"FE93",X"FE65",X"FE67",X"FEA3",X"FEF1",X"FF07",X"FF3E",X"FF6E",X"FF82",X"FFA0",X"FFD9",X"0000",X"FFD1",X"FFB4",X"FF9A",X"FF6E",
		X"FF55",X"FF43",X"FF7A",X"FF76",X"FF98",X"FFD0",X"FFFE",X"002C",X"0003",X"0000",X"0005",X"000D",X"0008",X"0030",X"001D",X"002F",
		X"0079",X"0067",X"0089",X"00DB",X"012E",X"016B",X"0149",X"0157",X"0160",X"0165",X"013A",X"0129",X"0119",X"00E8",X"00C5",X"00C8",
		X"00EC",X"00DF",X"00EE",X"0121",X"0115",X"00FC",X"013F",X"015D",X"0174",X"0156",X"0138",X"013B",X"010E",X"011E",X"0105",X"00CA",
		X"007B",X"004E",X"0038",X"0009",X"0002",X"FFD7",X"FFB8",X"FF91",X"FF81",X"FF7A",X"FF7E",X"FF70",X"FF4E",X"FF3C",X"FF0A",X"FED3",
		X"FE8C",X"FE49",X"FE10",X"FE1D",X"FE20",X"FE35",X"FE32",X"FE78",X"FE9D",X"FEB8",X"FEDE",X"FEF3",X"FEF3",X"FED0",X"FEBE",X"FECF",
		X"FEC8",X"FEE5",X"FF22",X"FF34",X"FF3E",X"FF64",X"FFA0",X"FFE0",X"0025",X"005A",X"0070",X"004D",X"0074",X"008C",X"008B",X"0092",
		X"00BB",X"00AE",X"0072",X"0062",X"0033",X"000C",X"FFFB",X"FFDB",X"FFDA",X"FFB2",X"FFE4",X"FFF4",X"FFF4",X"FFFF",X"000E",X"0007",
		X"0003",X"0014",X"0045",X"005D",X"0075",X"0089",X"0085",X"00BE",X"00FB",X"0153",X"0194",X"01CE",X"01B3",X"01AD",X"0175",X"013C",
		X"0122",X"00F4",X"00BD",X"009A",X"008A",X"00A2",X"00A5",X"00C0",X"0114",X"015D",X"01BA",X"01AF",X"01C9",X"01FF",X"01CB",X"01C8",
		X"01AE",X"018E",X"01B3",X"0186",X"0164",X"0152",X"0152",X"0147",X"00F8",X"00B8",X"0097",X"0085",X"0084",X"0055",X"0057",X"005A",
		X"0033",X"004F",X"006E",X"003F",X"001E",X"FFFD",X"FFCE",X"FFAD",X"FF8B",X"FF53",X"FF00",X"FECD",X"FF00",X"FF21",X"FF08",X"FEFD",
		X"FF11",X"FF0B",X"FEDC",X"FEBB",X"FEA2",X"FE6C",X"FE30",X"FDFC",X"FDEA",X"FE09",X"FE27",X"FE4A",X"FE61",X"FE96",X"FEC7",X"FED5",
		X"FED3",X"FEA7",X"FE8E",X"FE61",X"FE52",X"FE52",X"FE51",X"FE46",X"FE2B",X"FE51",X"FE53",X"FEA7",X"FED2",X"FF1B",X"FF2D",X"FF54",
		X"FF71",X"FF65",X"FF6B",X"FF43",X"FF0F",X"FEF3",X"FEFC",X"FEE0",X"FECB",X"FEF6",X"FF16",X"FEF7",X"FEDA",X"FEEF",X"FEE0",X"FECF",
		X"FEEA",X"FECF",X"FED2",X"FEE9",X"FF20",X"FF59",X"FF8E",X"FFC2",X"FFFB",X"0003",X"0001",X"0023",X"004D",X"0056",X"0043",X"0046",
		X"0068",X"006A",X"0094",X"00AA",X"0077",X"008B",X"0090",X"0075",X"006D",X"006C",X"0053",X"005C",X"007D",X"00BF",X"00BE",X"00DC",
		X"011E",X"0135",X"018A",X"01C4",X"01D8",X"01BC",X"0196",X"017C",X"0148",X"013B",X"012F",X"011A",X"010B",X"0124",X"0121",X"0118",
		X"0145",X"015E",X"0152",X"0150",X"018C",X"0172",X"0156",X"015A",X"016A",X"0169",X"014C",X"014F",X"0121",X"00F9",X"00E7",X"0107",
		X"0117",X"00F5",X"00C0",X"009B",X"008A",X"0077",X"0077",X"0033",X"FFF7",X"FFC3",X"FFDA",X"FFD2",X"FFC3",X"FFE6",X"FFF9",X"0010",
		X"0037",X"003D",X"0005",X"FFB3",X"FF79",X"FF25",X"FEF2",X"FED6",X"FEB4",X"FE8B",X"FE3F",X"FE47",X"FE78",X"FEC9",X"FEFC",X"FF37",
		X"FF4C",X"FF4C",X"FF6A",X"FF3A",X"FF0B",X"FEDB",X"FEB0",X"FE9C",X"FE75",X"FE84",X"FEB0",X"FED2",X"FEDA",X"FF0D",X"FF5E",X"FF68",
		X"FFA5",X"FFCA",X"FFC0",X"FF96",X"FF82",X"FFBB",X"FFAA",X"FF9D",X"FFCB",X"0000",X"FFEA",X"FFD5",X"FFF6",X"FFFF",X"FFBF",X"FFA6",
		X"FFCD",X"FFCD",X"FFD9",X"FFE8",X"002C",X"004B",X"007C",X"00BF",X"00A4",X"00A7",X"009F",X"0092",X"0087",X"0060",X"0073",X"0048",
		X"0068",X"006E",X"007B",X"0076",X"002F",X"0023",X"FFE6",X"000F",X"0026",X"0011",X"FFF4",X"FFED",X"001B",X"0030",X"0043",X"0053",
		X"001B",X"0012",X"001E",X"0029",X"0038",X"0032",X"0012",X"0000",X"FFFF",X"FFFE",X"0007",X"0023",X"FFF0",X"FFE0",X"0013",X"0044",
		X"0052",X"0036",X"0012",X"002A",X"0047",X"006E",X"0084",X"009E",X"00CB",X"00D0",X"00DA",X"00C7",X"00A8",X"00B2",X"00C2",X"00A8",
		X"00B0",X"00A4",X"00B9",X"00C3",X"00DE",X"0139",X"0156",X"0137",X"0130",X"00FE",X"00C6",X"0087",X"005B",X"FFFA",X"FFC6",X"FFB2",
		X"FFB6",X"FFA7",X"FFB0",X"FFDF",X"FFF6",X"003B",X"0089",X"0099",X"0096",X"008B",X"005E",X"007B",X"00A0",X"00AC",X"00B3",X"00B4",
		X"00A8",X"0092",X"0050",X"002D",X"0010",X"FFFE",X"FFF1",X"FFBC",X"FF84",X"FF6C",X"FF84",X"FF9C",X"FFB0",X"0007",X"001C",X"0027",
		X"0037",X"0049",X"0044",X"0048",X"0061",X"0065",X"002A",X"FFFB",X"FFEB",X"FFF0",X"FFEC",X"FFEC",X"FFD7",X"FFD6",X"FFE1",X"FFDD",
		X"FFC8",X"FFBA",X"FFBD",X"FFE7",X"FFD9",X"FFD6",X"FFA7",X"FF94",X"FF7B",X"FF6C",X"FF5C",X"FF58",X"FF76",X"FF7C",X"FF97",X"FFB7",
		X"0000",X"0013",X"003E",X"003D",X"005A",X"0048",X"005C",X"0069",X"0061",X"0047",X"0034",X"003B",X"003C",X"0049",X"0040",X"0058",
		X"0066",X"0069",X"0076",X"0093",X"0090",X"0070",X"005E",X"0059",X"0016",X"FFD2",X"FF6B",X"FEFF",X"FEDB",X"FED3",X"FEE7",X"FEEC",
		X"FF06",X"FF38",X"FF79",X"FFCD",X"0014",X"0040",X"0071",X"0081",X"00A3",X"00B5",X"00B2",X"00BC",X"00A4",X"00B6",X"00E6",X"0113",
		X"014D",X"0170",X"01CB",X"0205",X"021B",X"0250",X"0263",X"024C",X"021A",X"01DC",X"019E",X"017C",X"0143",X"0106",X"00D8",X"00BD",
		X"00B9",X"00A2",X"007D",X"0051",X"0030",X"FFE7",X"FF92",X"FF2B",X"FEBD",X"FE5A",X"FDF6",X"FDBE",X"FD6F",X"FD24",X"FCE4",X"FCE1",
		X"FCF9",X"FD43",X"FD70",X"FD8C",X"FDAB",X"FDD1",X"FE10",X"FE74",X"FEBC",X"FEE7",X"FEE1",X"FEE5",X"FEFA",X"FF05",X"FF33",X"FF50",
		X"FF74",X"FF8A",X"FFA6",X"FFEA",X"0035",X"00A5",X"00FD",X"0142",X"018B",X"01D1",X"020E",X"0255",X"029C",X"02B4",X"02D7",X"02D6",
		X"02FB",X"0326",X"0351",X"0341",X"034D",X"0352",X"0346",X"031B",X"0308",X"030C",X"02F6",X"02C9",X"0290",X"024F",X"01FC",X"01B2",
		X"0154",X"00B3",X"FFFF",X"FF31",X"FE4E",X"FD93",X"FCB0",X"FBDE",X"FAED",X"FA19",X"F997",X"F956",X"F943",X"F932",X"F918",X"F8F4",
		X"F90F",X"F935",X"F992",X"F9DA",X"FA1D",X"FA7B",X"FAE9",X"FB7C",X"FBFA",X"FC97",X"FD25",X"FDE6",X"FE78",X"FF0E",X"FFB8",X"0047",
		X"00AA",X"0104",X"014F",X"019A",X"01CA",X"01EA",X"0216",X"0242",X"027E",X"02B5",X"0307",X"0354",X"03BE",X"0457",X"04DC",X"0576",
		X"05E1",X"0637",X"069C",X"06F1",X"072F",X"0726",X"0714",X"06E9",X"06A3",X"064A",X"05E6",X"0574",X"0506",X"048C",X"0454",X"0403",
		X"0395",X"0324",X"02AE",X"0231",X"01A5",X"00EA",X"0014",X"FF48",X"FE66",X"FDA5",X"FCDA",X"FC26",X"FB9D",X"FB29",X"FAEC",X"FAAA",
		X"FA7C",X"FA59",X"FA51",X"FA42",X"FA36",X"FA41",X"FA23",X"FA2C",X"FA46",X"FA7B",X"FAC7",X"FB4B",X"FBEB",X"FC7C",X"FD0F",X"FDC7",
		X"FE70",X"FF09",X"FF96",X"0014",X"007B",X"00D0",X"0118",X"013D",X"0138",X"014F",X"016C",X"016A",X"016F",X"0166",X"0181",X"01A7",
		X"01BB",X"01E9",X"0202",X"0212",X"0217",X"0215",X"022B",X"0220",X"0205",X"01DA",X"01A7",X"0187",X"017B",X"0155",X"015A",X"014B",
		X"0167",X"017F",X"01A6",X"01F3",X"0211",X"022B",X"0236",X"0220",X"0208",X"01EC",X"01BA",X"0177",X"0122",X"00DA",X"00AB",X"0080",
		X"003D",X"0001",X"FFC2",X"FF72",X"FF03",X"FECB",X"FE89",X"FE23",X"FDC4",X"FD56",X"FCD1",X"FC60",X"FC0E",X"FBEE",X"FBCF",X"FBB6",
		X"FBA1",X"FBB2",X"FBD2",X"FC1C",X"FC94",X"FCE4",X"FD30",X"FD68",X"FD9E",X"FDDD",X"FE2C",X"FE59",X"FE8D",X"FEB2",X"FEDD",X"FF13",
		X"FF64",X"FFC9",X"0020",X"0067",X"009B",X"00C8",X"0104",X"0131",X"0147",X"0168",X"0153",X"0183",X"0198",X"01A7",X"01C1",X"0201",
		X"0257",X"02A1",X"02FF",X"033F",X"036C",X"0396",X"03C1",X"03F7",X"040F",X"0415",X"03F6",X"03F3",X"0414",X"041E",X"0439",X"0453",
		X"0483",X"049D",X"0485",X"0464",X"0451",X"0408",X"03AB",X"0341",X"02CA",X"0249",X"01B3",X"012E",X"00B1",X"004E",X"FFEC",X"FF9C",
		X"FF36",X"FEB8",X"FE5E",X"FE06",X"FD86",X"FCF4",X"FC4F",X"FBAE",X"FB30",X"FAA6",X"FA2E",X"F9B3",X"F940",X"F8EA",X"F8C2",X"F8D0",
		X"F8CD",X"F8CC",X"F8E9",X"F92B",X"F9A9",X"FA29",X"FA96",X"FB10",X"FB8B",X"FBF8",X"FC66",X"FCC3",X"FD3C",X"FDC7",X"FE4E",X"FEB3",
		X"FF13",X"FF89",X"001E",X"00B5",X"0118",X"017E",X"01B9",X"01B0",X"01C9",X"01D2",X"01C9",X"0198",X"014A",X"0107",X"00FE",X"0109",
		X"0142",X"017B",X"01C3",X"0239",X"02C4",X"033E",X"03A8",X"0400",X"0434",X"0446",X"0451",X"045E",X"045F",X"0447",X"0429",X"0446",
		X"0466",X"049F",X"04DD",X"04EC",X"04DF",X"04F0",X"04C6",X"0467",X"03F3",X"034F",X"027A",X"01C7",X"010F",X"0043",X"FF8F",X"FF04",
		X"FE94",X"FE41",X"FE27",X"FE06",X"FDE2",X"FDEA",X"FE1C",X"FE3B",X"FE56",X"FE8E",X"FEB9",X"FEC3",X"FEED",X"FF14",X"FF4E",X"FF73",
		X"FFA1",X"FFF2",X"0026",X"0097",X"00F0",X"0121",X"016A",X"01AD",X"01A3",X"0179",X"012A",X"00C9",X"0045",X"FFA0",X"FEFF",X"FE40",
		X"FD90",X"FCEB",X"FC7D",X"FC29",X"FBEE",X"FBDD",X"FBFC",X"FC28",X"FC39",X"FC55",X"FC88",X"FCB0",X"FCE2",X"FD19",X"FD4A",X"FD7C",
		X"FDBD",X"FE0E",X"FE5E",X"FECB",X"FF3D",X"FF88",X"FFEC",X"0041",X"0086",X"00B2",X"00E2",X"00F6",X"00E4",X"00C0",X"0094",X"0078",
		X"0045",X"0017",X"FFBB",X"FF6D",X"FF18",X"FEBE",X"FE5F",X"FE0D",X"FDD6",X"FDBE",X"FD9F",X"FDA3",X"FDBF",X"FE02",X"FE1B",X"FE28",
		X"FE4E",X"FE6D",X"FE85",X"FE71",X"FE5D",X"FE39",X"FE2E",X"FE32",X"FE1C",X"FDEF",X"FDD8",X"FDF0",X"FDF5",X"FE01",X"FE17",X"FE3E",
		X"FE5D",X"FE5D",X"FE68",X"FE96",X"FECC",X"FF22",X"FFB0",X"0006",X"005A",X"00B3",X"0127",X"01BE",X"023A",X"02CB",X"0336",X"0389",
		X"03ED",X"0444",X"04A1",X"0513",X"0562",X"058B",X"05DD",X"0626",X"067E",X"06D5",X"073A",X"078C",X"07C9",X"0817",X"0842",X"085C",
		X"0856",X"081C",X"07F4",X"07A5",X"074A",X"06E3",X"0688",X"0661",X"062E",X"05EA",X"05B4",X"0579",X"0556",X"053A",X"04F8",X"0472",
		X"03B7",X"0301",X"0235",X"0174",X"009E",X"FFC7",X"FEF7",X"FE2F",X"FD93",X"FD31",X"FD0D",X"FCF8",X"FCDE",X"FCEC",X"FD12",X"FD0B",
		X"FD0B",X"FCDD",X"FC95",X"FC55",X"FBF7",X"FBA6",X"FB42",X"FAFA",X"FAD1",X"FADF",X"FAF3",X"FB26",X"FB6D",X"FBA2",X"FBE8",X"FC41",
		X"FC80",X"FC9A",X"FCA9",X"FCA4",X"FC9C",X"FC95",X"FC9D",X"FCA6",X"FC95",X"FCAA",X"FCC6",X"FCCB",X"FCD7",X"FD04",X"FD22",X"FD19",
		X"FD0D",X"FCFD",X"FCD6",X"FC91",X"FC58",X"FC26",X"FBE3",X"FBB2",X"FB64",X"FAF3",X"FA98",X"FA2D",X"F9E4",X"F9B0",X"F998",X"F989",
		X"F9AE",X"F9EF",X"FA5D",X"FAB8",X"FB08",X"FB3C",X"FB6B",X"FBC4",X"FBE6",X"FC03",X"FC03",X"FC20",X"FC79",X"FCEA",X"FD80",X"FE27",
		X"FEBB",X"FF59",X"0003",X"00A3",X"0106",X"0161",X"018F",X"019B",X"01CF",X"01ED",X"0206",X"0235",X"0275",X"02D1",X"033D",X"03AB",
		X"044A",X"04E4",X"0586",X"063C",X"06C5",X"073C",X"0780",X"07B5",X"07F7",X"07E9",X"07C9",X"0791",X"0768",X"072A",X"06D5",X"069F",
		X"067D",X"0637",X"05F3",X"05B2",X"0551",X"04E8",X"046A",X"03B5",X"0326",X"02AD",X"0240",X"01B7",X"013B",X"00CE",X"0056",X"0045",
		X"0030",X"0026",X"0023",X"0026",X"0040",X"006F",X"00A9",X"00E7",X"0102",X"013B",X"0175",X"01CF",X"024B",X"028F",X"0311",X"0379",
		X"03D8",X"0443",X"0496",X"0500",X"052D",X"052C",X"0530",X"04FB",X"04D3",X"04B5",X"04B5",X"04AE",X"045A",X"0438",X"03E7",X"0392",
		X"0357",X"030F",X"02BA",X"0257",X"01D3",X"013D",X"00CC",X"0057",X"0001",X"FF73",X"FEBF",X"FE1F",X"FD8D",X"FD28",X"FCC8",X"FC5A",
		X"FBDE",X"FB5F",X"FAE1",X"FA83",X"FA13",X"F9C5",X"F950",X"F8C1",X"F86A",X"F81A",X"F7AD",X"F730",X"F68C",X"F5DF",X"F524",X"F46C",
		X"F3CC",X"F33C",X"F2D2",X"F297",X"F26F",X"F279",X"F2AD",X"F31D",X"F3CB",X"F45E",X"F4FD",X"F59B",X"F65E",X"F741",X"F807",X"F8B5",
		X"F97B",X"FA45",X"FB0B",X"FBD7",X"FCC0",X"FDC0",X"FEBB",X"FFAC",X"0086",X"0161",X"0226",X"02BC",X"032D",X"03B7",X"041E",X"046F",
		X"04C5",X"051E",X"0576",X"05C8",X"0631",X"0687",X"06DB",X"06FB",X"0705",X"070A",X"0702",X"06CD",X"0682",X"063D",X"0619",X"05F9",
		X"05DF",X"05DA",X"05F5",X"0632",X"0656",X"069E",X"06E8",X"072C",X"073F",X"071A",X"06F4",X"06BB",X"065F",X"0618",X"05CB",X"0578",
		X"0542",X"04FA",X"04AC",X"0462",X"0435",X"03FC",X"03AB",X"0361",X"0339",X"033F",X"0356",X"0372",X"039B",X"03D3",X"0417",X"0456",
		X"04A5",X"04CA",X"04D1",X"04D0",X"049D",X"0444",X"03D1",X"0358",X"02D5",X"025E",X"0200",X"0178",X"00EA",X"0091",X"0031",X"FFC4",
		X"FF84",X"FF47",X"FF0F",X"FEB9",X"FE62",X"FE0B",X"FDA3",X"FD64",X"FD14",X"FC9E",X"FC48",X"FBE0",X"FB90",X"FB61",X"FB40",X"FB10",
		X"FADC",X"FAB4",X"FA69",X"FA4E",X"FA4B",X"FA31",X"F9FC",X"F9DF",X"F9AB",X"F999",X"F992",X"F9A9",X"F9C1",X"F9E3",X"FA16",X"FA3B",
		X"FA34",X"FA16",X"F9FC",X"F9CE",X"F977",X"F951",X"F925",X"F90B",X"F901",X"F90B",X"F944",X"F99F",X"FA0C",X"FA7C",X"FAF3",X"FB6E",
		X"FBFA",X"FC75",X"FCF1",X"FD33",X"FD88",X"FDD3",X"FE0C",X"FE60",X"FEC7",X"FF06",X"FF4C",X"FF7B",X"FF9E",X"FF9D",X"FF9A",X"FF8D",
		X"FF8C",X"FFB0",X"FFC4",X"FFF2",X"003C",X"0091",X"00E2",X"0153",X"01B1",X"021E",X"0268",X"02A3",X"02DD",X"02ED",X"0300",X"031C",
		X"0313",X"031A",X"0321",X"033D",X"0360",X"03A1",X"0417",X"0486",X"0513",X"057F",X"05EB",X"0648",X"06AB",X"06EB",X"0725",X"075C",
		X"078F",X"079A",X"07B6",X"07E2",X"0810",X"0822",X"0806",X"07F2",X"07E1",X"07E4",X"07CA",X"0772",X"0717",X"06BE",X"0677",X"0662",
		X"066B",X"067D",X"0646",X"0601",X"05A2",X"051A",X"047E",X"03C3",X"02D7",X"01C1",X"00B1",X"FFA5",X"FEE8",X"FE4F",X"FDA7",X"FD3E",
		X"FCE5",X"FCBE",X"FCBC",X"FCD8",X"FD06",X"FD1C",X"FCF0",X"FCA1",X"FC65",X"FC05",X"FBA5",X"FB2D",X"FAAE",X"FA43",X"F9E6",X"F9AA",
		X"F9A5",X"F9CC",X"F9E3",X"F9FE",X"FA33",X"FA83",X"FAE0",X"FB39",X"FBA2",X"FBB1",X"FBAD",X"FBC9",X"FBCB",X"FBD6",X"FBE3",X"FBCC",
		X"FB9D",X"FB66",X"FB58",X"FB76",X"FB8F",X"FBCD",X"FBF3",X"FC23",X"FC6A",X"FCC4",X"FD39",X"FD7F",X"FDC4",X"FDF8",X"FE37",X"FE6C",
		X"FEBB",X"FF0C",X"FF3A",X"FF55",X"FF6C",X"FF65",X"FF82",X"FFC1",X"FFF8",X"0037",X"0048",X"0073",X"00B2",X"00EC",X"0155",X"01A6",
		X"01C4",X"01A1",X"015F",X"013A",X"0106",X"00DC",X"00CC",X"00A8",X"008F",X"0065",X"0029",X"FFF2",X"FFBD",X"FF60",X"FEF1",X"FE75",
		X"FE07",X"FDBC",X"FDB9",X"FDCD",X"FDCA",X"FE05",X"FE76",X"FEF4",X"FFA3",X"0059",X"00D9",X"0153",X"01AC",X"01EA",X"021E",X"0263",
		X"02C1",X"02F1",X"0330",X"0354",X"03B2",X"042C",X"048F",X"0539",X"05E5",X"0678",X"06CA",X"0711",X"0750",X"0768",X"073B",X"070E",
		X"06E4",X"06D8",X"06B9",X"06BD",X"06C0",X"06B3",X"068D",X"0662",X"060D",X"05B9",X"0538",X"04C0",X"045A",X"03FB",X"03B6",X"038A",
		X"0385",X"038F",X"03A1",X"03B0",X"03AA",X"036C",X"0314",X"02AE",X"0211",X"0139",X"006D",X"FFA4",X"FEF4",X"FE16",X"FD66",X"FCDA",
		X"FC2F",X"FBA7",X"FB39",X"FACD",X"FA6B",X"F9FD",X"F996",X"F948",X"F8DB",X"F87A",X"F806",X"F796",X"F73A",X"F70B",X"F6F9",X"F6DC",
		X"F6B9",X"F6A8",X"F69F",X"F697",X"F6A1",X"F694",X"F68B",X"F68D",X"F6C2",X"F6CA",X"F6F5",X"F71F",X"F77D",X"F7CD",X"F832",X"F8F8",
		X"F999",X"FA33",X"FAB1",X"FB23",X"FBA7",X"FC40",X"FCBD",X"FD2E",X"FD69",X"FDD8",X"FE3E",X"FEAD",X"FF33",X"FFB4",X"006C",X"010C",
		X"018F",X"021D",X"029E",X"031B",X"0371",X"03C6",X"03FD",X"0417",X"045D",X"04C0",X"053D",X"05C3",X"064E",X"06CC",X"073D",X"0783",
		X"07DB",X"07F2",X"07F9",X"07F5",X"07D0",X"07B4",X"07B7",X"07C5",X"07D9",X"07FB",X"0818",X"0824",X"0827",X"083E",X"082B",X"080A",
		X"07AC",X"0742",X"06E8",X"068C",X"0624",X"05AF",X"0552",X"050F",X"04D7",X"04C2",X"04A8",X"049C",X"0478",X"042F",X"03D3",X"033A",
		X"02AD",X"0229",X"01A0",X"0117",X"0097",X"0024",X"FFD1",X"FF70",X"FF31",X"FED3",X"FE4B",X"FDBE",X"FCFF",X"FC1F",X"FB3E",X"FA6C",
		X"F9C6",X"F950",X"F913",X"F90A",X"F93D",X"F998",X"FA26",X"FAD5",X"FB64",X"FBC8",X"FC11",X"FC6E",X"FCE3",X"FD64",X"FDB1",X"FDDE",
		X"FE0E",X"FE23",X"FE38",X"FE47",X"FE39",X"FE1E",X"FDD7",X"FD95",X"FD77",X"FD5F",X"FD71",X"FD83",X"FDA7",X"FDA5",X"FDB7",X"FDDF",
		X"FE12",X"FE30",X"FE37",X"FE3F",X"FE4C",X"FE62",X"FE65",X"FE67",X"FE62",X"FE68",X"FE6C",X"FE84",X"FE8B",X"FEA2",X"FEBD",X"FED8",
		X"FEC6",X"FEA6",X"FE57",X"FE06",X"FDC4",X"FD3A",X"FC97",X"FBEA",X"FB3B",X"FA98",X"FA38",X"F9FB",X"FA03",X"FA1A",X"FA5A",X"FABF",
		X"FB59",X"FC37",X"FCD7",X"FD70",X"FDF0",X"FE50",X"FE84",X"FEBC",X"FEDE",X"FEFC",X"FEF3",X"FEF6",X"FF37",X"FFA2",X"002C",X"00E2",
		X"01AA",X"0275",X"0326",X"03A1",X"03FD",X"042F",X"042D",X"0425",X"0433",X"0462",X"049F",X"04F8",X"0594",X"0630",X"06D0",X"07AC",
		X"0887",X"0973",X"0A31",X"0ACA",X"0B28",X"0B25",X"0B14",X"0ADF",X"0A9D",X"0A3A",X"09F4",X"099F",X"0930",X"08D6",X"089A",X"083A",
		X"07EF",X"0783",X"06E2",X"0646",X"0562",X"046D",X"0357",X"0229",X"00EF",X"FFD4",X"FEDC",X"FE1F",X"FD93",X"FD08",X"FC81",X"FBF4",
		X"FB8D",X"FB1E",X"FA97",X"F9EB",X"F935",X"F873",X"F7F1",X"F765",X"F6E2",X"F67B",X"F615",X"F5D1",X"F5B6",X"F5D3",X"F5EB",X"F61D",
		X"F661",X"F6B5",X"F73C",X"F7E6",X"F888",X"F941",X"FA09",X"FAD7",X"FB8A",X"FC18",X"FC97",X"FCF6",X"FD39",X"FD75",X"FD90",X"FD94",
		X"FD9D",X"FDD4",X"FE16",X"FE7D",X"FEB9",X"FF09",X"FF92",X"002D",X"00C6",X"0143",X"0198",X"01D9",X"020A",X"0232",X"025B",X"0262",
		X"0273",X"0279",X"0293",X"02B6",X"02D7",X"02E7",X"02FB",X"030F",X"0305",X"02FA",X"0327",X"02F3",X"02DC",X"02CE",X"028D",X"024E",
		X"01F9",X"01C1",X"01A8",X"0193",X"01A3",X"01C8",X"01F0",X"023B",X"0262",X"0251",X"0232",X"020A",X"01D1",X"017E",X"00FF",X"0095",
		X"004C",X"FFE8",X"FFC9",X"FFC4",X"FFBF",X"FFE8",X"0057",X"00A2",X"00D9",X"012C",X"0161",X"018A",X"017C",X"0152",X"0127",X"0106",
		X"00EB",X"00C2",X"0097",X"007A",X"0087",X"008F",X"00B2",X"00CF",X"0106",X"0136",X"0126",X"0100",X"00B1",X"007A",X"0028",X"FFE1",
		X"FF82",X"FF1E",X"FECB",X"FE7D",X"FE59",X"FE48",X"FE3A",X"FE32",X"FE52",X"FE5C",X"FE80",X"FEBB",X"FEB8",X"FEB9",X"FED1",X"FEF1",
		X"FF0F",X"FF36",X"FF8C",X"FFC7",X"FFD4",X"0008",X"005F",X"00C4",X"00E5",X"00F5",X"00DF",X"00BB",X"00AD",X"00B3",X"008D",X"0072",
		X"004A",X"0039",X"0043",X"0033",X"005E",X"006A",X"004F",X"003F",X"003F",X"006A",X"00A0",X"00ED",X"012D",X"015E",X"0199",X"01D0",
		X"0211",X"0216",X"021F",X"0221",X"01B7",X"0139",X"00D5",X"0069",X"0014",X"FFB4",X"FF65",X"FF45",X"FF38",X"FF42",X"FF5A",X"FF55",
		X"FF47",X"FF34",X"FF19",X"FEC1",X"FE87",X"FE31",X"FDB8",X"FD2F",X"FCD4",X"FCA4",X"FC80",X"FC9B",X"FCCB",X"FD1B",X"FD80",X"FE03",
		X"FE86",X"FEEF",X"FF41",X"FFBF",X"001B",X"0055",X"005F",X"0073",X"009F",X"00A3",X"00CB",X"00ED",X"00FC",X"012F",X"0161",X"01C1",
		X"0219",X"0256",X"0284",X"0291",X"02A2",X"0287",X"026A",X"025D",X"024D",X"023E",X"0230",X"0218",X"01E9",X"01D4",X"01C8",X"01D5",
		X"01BF",X"01C8",X"01C4",X"01B7",X"01B5",X"01AC",X"01A6",X"0183",X"0159",X"0139",X"0142",X"012E",X"011C",X"00F3",X"00C9",X"006A",
		X"FFE9",X"FF72",X"FF21",X"FEC3",X"FE27",X"FDA8",X"FD3E",X"FCB2",X"FC27",X"FB8B",X"FAC6",X"F9EF",X"F91A",X"F864",X"F77C",X"F6D8",
		X"F672",X"F630",X"F612",X"F63A",X"F6AC",X"F737",X"F7E7",X"F896",X"F944",X"F9D5",X"FA5B",X"FAE2",X"FB51",X"FBCB",X"FC45",X"FCB0",
		X"FD2D",X"FDCE",X"FE84",X"FF4B",X"000D",X"00C7",X"0175",X"0217",X"02CC",X"0350",X"03C2",X"03FF",X"0420",X"043B",X"0454",X"04A2",
		X"04B7",X"04C7",X"04EB",X"0525",X"0590",X"0601",X"06B4",X"073E",X"07D7",X"085F",X"08E3",X"0943",X"099F",X"09C5",X"09AC",X"0972",
		X"0955",X"0920",X"08E3",X"08B8",X"0867",X"07FA",X"076B",X"06EE",X"065C",X"0596",X"04C4",X"03BF",X"0279",X"0156",X"004D",X"FF7A",
		X"FE87",X"FDE5",X"FD57",X"FCE1",X"FCAA",X"FCC1",X"FD1B",X"FD66",X"FDAC",X"FDDD",X"FE18",X"FE4B",X"FE94",X"FE9F",X"FEAD",X"FE9B",
		X"FE6E",X"FE43",X"FE1A",X"FE2A",X"FE15",X"FDCD",X"FD7C",X"FD4A",X"FD26",X"FD28",X"FD20",X"FD21",X"FD18",X"FD0F",X"FD40",X"FD79",
		X"FDB8",X"FDE9",X"FE22",X"FE4D",X"FE60",X"FE73",X"FE8B",X"FEA6",X"FE9A",X"FEB4",X"FEDC",X"FEFB",X"FF36",X"FF68",X"FFA0",X"FFCB",
		X"FFE6",X"FFE1",X"FFBD",X"FF87",X"FF55",X"FF1B",X"FECF",X"FE48",X"FDBB",X"FD2A",X"FC7A",X"FBAE",X"FB05",X"FA76",X"FA0A",X"F9D7",
		X"F9BE",X"F9C6",X"F9F0",X"FA66",X"FAE4",X"FB83",X"FC13",X"FC67",X"FC9C",X"FCA9",X"FCA3",X"FC72",X"FC14",X"FBB8",X"FB90",X"FB91",
		X"FBBA",X"FC32",X"FCCB",X"FD5C",X"FE40",X"FF22",X"0002",X"00D8",X"01A5",X"021E",X"0257",X"0260",X"023C",X"021B",X"020E",X"020B",
		X"01F3",X"0220",X"02A8",X"0360",X"040B",X"04BF",X"0578",X"061C",X"067F",X"0698",X"068E",X"0673",X"0636",X"05C7",X"053C",X"04C1",
		X"0466",X"0459",X"0434",X"0448",X"0453",X"043D",X"0456",X"0485",X"04BE",X"04F1",X"0523",X"051A",X"04F5",X"04F3",X"04C3",X"049B",
		X"0477",X"0452",X"0409",X"03BC",X"0369",X"0315",X"02E6",X"029B",X"023D",X"01CB",X"0164",X"00E5",X"0077",X"FFF4",X"FF5C",X"FEB9",
		X"FE52",X"FDCF",X"FD6A",X"FD49",X"FD5B",X"FD92",X"FDCB",X"FE2F",X"FE94",X"FEF0",X"FF5E",X"FFB6",X"FFEA",X"FFDD",X"FFA8",X"FF60",
		X"FEF9",X"FE72",X"FDC3",X"FCE8",X"FC17",X"FB2E",X"FA5F",X"F9BA",X"F925",X"F8C4",X"F88F",X"F889",X"F8C1",X"F909",X"F960",X"F9A6",
		X"F9E9",X"FA2D",X"FA68",X"FAA5",X"FA9B",X"FAA7",X"FACF",X"FB12",X"FB88",X"FC02",X"FCAE",X"FD7A",X"FE54",X"FF35",X"FFF0",X"00B0",
		X"013D",X"01A7",X"0225",X"0284",X"029E",X"0291",X"0242",X"01FC",X"01F1",X"0214",X"0262",X"02BD",X"0346",X"03C7",X"043C",X"04F1",
		X"05A5",X"064F",X"06C2",X"06F5",X"0716",X"0721",X"0759",X"07C8",X"0813",X"083A",X"083B",X"082A",X"081D",X"07FE",X"07E3",X"0773",
		X"06BF",X"05F6",X"052B",X"045B",X"0360",X"0275",X"0182",X"0097",X"FF9E",X"FE96",X"FDD5",X"FD0D",X"FC3B",X"FB89",X"FAD1",X"FA5B",
		X"FA0E",X"F9E2",X"F9EB",X"FA26",X"FA56",X"FAAD",X"FB15",X"FB69",X"FB97",X"FB98",X"FBAB",X"FB98",X"FB74",X"FB64",X"FB6C",X"FB84",
		X"FB7D",X"FB81",X"FBB2",X"FBC2",X"FBC8",X"FBD4",X"FBB6",X"FB91",X"FB69",X"FB21",X"FADB",X"FAC3",X"FABE",X"FABD",X"FAE7",X"FB55",
		X"FBE0",X"FC58",X"FCEB",X"FD62",X"FDBC",X"FE1F",X"FE79",X"FEB1",X"FEBF",X"FEB2",X"FEBC",X"FED3",X"FF14",X"FF3E",X"FF77",X"FFA7",
		X"FFC5",X"FFF7",X"0020",X"0072",X"00A7",X"00DD",X"00F3",X"010A",X"0148",X"018F",X"01BF",X"01E5",X"022F",X"0263",X"025F",X"027C",
		X"0282",X"024F",X"0216",X"01BA",X"015C",X"0111",X"00DD",X"00B0",X"0098",X"00C1",X"0103",X"0177",X"0201",X"02AA",X"0345",X"03BE",
		X"042E",X"0476",X"04C1",X"04DB",X"04C1",X"049B",X"0455",X"042E",X"0428",X"0401",X"03EB",X"0406",X"0439",X"044B",X"0434",X"0447",
		X"044E",X"0413",X"03D7",X"0398",X"0366",X"0341",X"0312",X"02E1",X"02BE",X"02BD",X"02B3",X"026C",X"0238",X"0207",X"01B2",X"0139",
		X"00D2",X"005E",X"0010",X"FFF6",X"FFE1",X"FFE2",X"0010",X"0081",X"0119",X"01D2",X"0278",X"0319",X"038D",X"03EA",X"040E",X"0411",
		X"03F6",X"0399",X"031B",X"0296",X"0234",X"01AE",X"0153",X"00F7",X"008D",X"0047",X"0006",X"FFE5",X"FF9E",X"FF51",X"FEEC",X"FE84",
		X"FE18",X"FDE2",X"FD9F",X"FD56",X"FCFC",X"FC99",X"FC27",X"FBBB",X"FB3D",X"FA94",X"F9C9",X"F8EE",X"F82A",X"F77D",X"F716",X"F6BA",
		X"F699",X"F6C0",X"F704",X"F741",X"F7BF",X"F850",X"F8D3",X"F927",X"F972",X"F9C2",X"F9D1",X"FA04",X"FA37",X"FA6A",X"FACB",X"FB13",
		X"FB71",X"FBDD",X"FC43",X"FCBF",X"FD43",X"FD9A",X"FDF5",X"FE1F",X"FE50",X"FE45",X"FE2F",X"FE2F",X"FE27",X"FE3E",X"FE72",X"FEC7",
		X"FF15",X"FF90",X"0046",X"00F2",X"01AF",X"026A",X"02F6",X"03A0",X"0444",X"04DB",X"0559",X"05C2",X"05FE",X"0602",X"05F5",X"05F5",
		X"05FB",X"05DC",X"05CD",X"05C7",X"05AE",X"05B1",X"05CB",X"060A",X"0633",X"061F",X"05FC",X"05BA",X"055C",X"04F4",X"047C",X"03F1",
		X"0329",X"027D",X"01DC",X"0188",X"0161",X"0148",X"0162",X"0146",X"0142",X"015F",X"017D",X"01B3",X"01CC",X"01D3",X"01BD",X"01AD",
		X"01AF",X"01CF",X"01D9",X"01D6",X"01AC",X"014A",X"0102",X"00DB",X"00B3",X"006E",X"0030",X"FFC8",X"FF42",X"FEC7",X"FE3A",X"FDC2",
		X"FD20",X"FC80",X"FC0E",X"FBA7",X"FB68",X"FB75",X"FBBE",X"FC3A",X"FC98",X"FCF3",X"FD3E",X"FD9C",X"FDF2",X"FDE0",X"FDBB",X"FD81",
		X"FD42",X"FD10",X"FCDC",X"FCD4",X"FCEF",X"FD3F",X"FDCE",X"FE76",X"FF55",X"002D",X"012A",X"01F7",X"0266",X"029A",X"02B9",X"02E0",
		X"02B9",X"0273",X"020A",X"01B5",X"0168",X"0128",X"00E7",X"0082",X"006F",X"003D",X"001B",X"FFDB",X"FFC3",X"FFA7",X"FFB3",X"FFCB",
		X"FFE6",X"001B",X"0070",X"00C8",X"011B",X"018A",X"01EA",X"0218",X"0205",X"01CC",X"0166",X"00EC",X"0068",X"FFF3",X"FF70",X"FEEB",
		X"FE4F",X"FDA9",X"FD15",X"FCA5",X"FC31",X"FBA7",X"FB22",X"FAB9",X"FA3E",X"FA12",X"F9E8",X"F9BC",X"F98D",X"F96F",X"F983",X"F98C",
		X"F9C7",X"FA1D",X"FA44",X"FA72",X"FAA7",X"FB1A",X"FBA5",X"FC24",X"FCB1",X"FD6A",X"FE37",X"FF00",X"FFD8",X"00A5",X"015A",X"01C8",
		X"020D",X"01E4",X"01A2",X"0149",X"00D0",X"006E",X"0011",X"FFDE",X"FFDB",X"FFED",X"005E",X"00FB",X"01C2",X"0286",X"0336",X"03DC",
		X"046F",X"050C",X"057A",X"05BE",X"05D7",X"05C4",X"05B3",X"057E",X"055B",X"0561",X"0547",X"054E",X"0565",X"059B",X"05E8",X"0622",
		X"068F",X"06D0",X"0703",X"0735",X"0744",X"0755",X"0751",X"0767",X"0784",X"07C5",X"07FC",X"0845",X"087B",X"08B6",X"0902",X"0903",
		X"08F0",X"08A0",X"084B",X"07B3",X"070B",X"0690",X"0602",X"0557",X"04D1",X"0488",X"0426",X"03DE",X"0364",X"0312",X"029D",X"01D5",
		X"010B",X"0008",X"FEC3",X"FD65",X"FC05",X"FAA8",X"F987",X"F876",X"F7C3",X"F727",X"F6E1",X"F6DB",X"F6EC",X"F71D",X"F76F",X"F7DE",
		X"F823",X"F85B",X"F875",X"F84A",X"F81D",X"F7F3",X"F7A8",X"F756",X"F6F2",X"F6A9",X"F689",X"F6AC",X"F6E2",X"F729",X"F7A9",X"F7FB",
		X"F84C",X"F8CA",X"F931",X"F95D",X"F951",X"F95E",X"F960",X"F9AB",X"FA00",X"FA56",X"FAB1",X"FB2E",X"FBD2",X"FC80",X"FCF0",X"FD6B",
		X"FDD6",X"FE0E",X"FE47",X"FE7F",X"FECA",X"FEC6",X"FEDE",X"FEC9",X"FE86",X"FE3F",X"FE10",X"FDCD",X"FDA3",X"FD75",X"FD2A",X"FD02",
		X"FCE7",X"FCCE",X"FCB5",X"FC9C",X"FC5D",X"FC13",X"FBE6",X"FBDD",X"FC1F",X"FC61",X"FC8B",X"FC9F",X"FCF9",X"FD63",X"FDD3",X"FE61",
		X"FEEB",X"FF57",X"FFD2",X"0074",X"0129",X"01EE",X"02C0",X"0386",X"0436",X"04F5",X"05CD",X"06A0",X"0765",X"0836",X"08E6",X"0979",
		X"0A05",X"0A78",X"0AF4",X"0B77",X"0BCE",X"0C05",X"0C29",X"0C32",X"0C11",X"0BF8",X"0BBD",X"0B46",X"0ADF",X"0A74",X"0A34",X"0A18",
		X"0A04",X"0A13",X"0A3B",X"0A86",X"0AD1",X"0AD4",X"0AD4",X"0AB8",X"0A63",X"0A06",X"0955",X"089D",X"07C6",X"0714",X"066F",X"05DA",
		X"0521",X"049C",X"0446",X"03D3",X"0362",X"02D3",X"0242",X"01A2",X"0112",X"0035",X"FF68",X"FE9A",X"FDC3",X"FCFA",X"FC3E",X"FB7E",
		X"FAC0",X"F9FB",X"F954",X"F8D1",X"F850",X"F7DE",X"F780",X"F746",X"F6FF",X"F6EE",X"F6F6",X"F71D",X"F74F",X"F7A3",X"F7EB",X"F7F5",
		X"F7DB",X"F7AF",X"F75C",X"F6FD",X"F686",X"F5EB",X"F533",X"F47C",X"F40A",X"F3CD",X"F3B5",X"F3A6",X"F3BE",X"F417",X"F495",X"F519",
		X"F5B5",X"F662",X"F6CA",X"F720",X"F758",X"F776",X"F789",X"F7AB",X"F7CE",X"F831",X"F8D8",X"F9AC",X"FAAB",X"FBD2",X"FD09",X"FE3A",
		X"FF82",X"008C",X"0178",X"0228",X"029A",X"02E2",X"0327",X"0331",X"0331",X"0348",X"0366",X"039F",X"03E9",X"044E",X"04A4",X"051E",
		X"05AA",X"0642",X"06ED",X"0775",X"0802",X"0868",X"08D1",X"092D",X"0974",X"09A2",X"09AC",X"09C3",X"09E5",X"09E4",X"09D8",X"09AD",
		X"0967",X"0934",X"08E0",X"0880",X"07F9",X"0778",X"0723",X"06DB",X"0671",X"05EA",X"0566",X"04D0",X"0461",X"03E0",X"038A",X"0319",
		X"02BD",X"028E",X"026B",X"0254",X"0271",X"0270",X"0270",X"0289",X"0276",X"0288",X"0267",X"025A",X"0220",X"0202",X"01E4",X"01D8",
		X"01A4",X"016F",X"0147",X"0127",X"0116",X"0118",X"0131",X"0132",X"0124",X"00EE",X"009E",X"004C",X"0011",X"FFBE",X"FF41",X"FED2",
		X"FE43",X"FDA1",X"FD2B",X"FCFD",X"FCDC",X"FCCD",X"FCAE",X"FC83",X"FC28",X"FB9E",X"FB28",X"FA5C",X"F97E",X"F88D",X"F778",X"F660",
		X"F569",X"F4C0",X"F439",X"F3D7",X"F3AD",X"F3C2",X"F3ED",X"F450",X"F4DC",X"F58E",X"F61C",X"F68C",X"F72C",X"F7D8",X"F882",X"F924",
		X"F9AE",X"FA35",X"FAC2",X"FB48",X"FBDB",X"FC49",X"FCAC",X"FD1D",X"FD7D",X"FDEE",X"FE62",X"FED5",X"FF35",X"FF71",X"FFA1",X"FFA7",
		X"FFC7",X"FFA9",X"FF8B",X"FF28",X"FEF2",X"FEB9",X"FE78",X"FE83",X"FE8A",X"FEC5",X"FF2C",X"FFD6",X"00A6",X"0174",X"024E",X"0330",
		X"041E",X"04DA",X"0583",X"0626",X"06B6",X"0700",X"0724",X"072B",X"072A",X"0739",X"0735",X"0733",X"0716",X"06FE",X"06F2",X"06E1",
		X"06D2",X"06BC",X"0696",X"0654",X"061D",X"05D9",X"0594",X"0564",X"0526",X"050A",X"04E8",X"04FC",X"052B",X"05A4",X"05F3",X"063B",
		X"069C",X"06D2",X"06F0",X"06F2",X"06D9",X"06A5",X"0644",X"05D8",X"0560",X"04D8",X"045E",X"041A",X"03BD",X"0386",X"0367",X"033B",
		X"0309",X"02BE",X"0283",X"0225",X"01A4",X"0110",X"0067",X"FFB7",X"FF07",X"FE59",X"FDBE",X"FD34",X"FCB3",X"FC42",X"FBF9",X"FBAD",
		X"FB7B",X"FB46",X"FB0A",X"FA9D",X"FA2C",X"F9AD",X"F959",X"F8E4",X"F890",X"F852",X"F81B",X"F80F",X"F822",X"F876",X"F8AA",X"F8DC",
		X"F928",X"F993",X"F9E4",X"FA29",X"FA74",X"FADC",X"FB1C",X"FB38",X"FB5F",X"FB6F",X"FB9A",X"FBAA",X"FBD9",X"FC13",X"FC35",X"FC84",
		X"FCE1",X"FD5E",X"FDEF",X"FE6D",X"FED6",X"FF51",X"FFDF",X"0044",X"00B1",X"011A",X"014E",X"0187",X"01B1",X"01FC",X"024A",X"02AC",
		X"02FC",X"035B",X"038C",X"03CA",X"040B",X"040D",X"0404",X"03C9",X"03A0",X"033A",X"02C9",X"026E",X"020E",X"019D",X"0145",X"0123",
		X"011C",X"0129",X"014A",X"0145",X"0132",X"0122",X"011B",X"0120",X"0122",X"0141",X"0144",X"0134",X"0141",X"017C",X"01D3",X"0244",
		X"02BB",X"032F",X"038D",X"03C7",X"0415",X"045A",X"048D",X"0486",X"0484",X"0472",X"0446",X"0412",X"03D4",X"038B",X"032F",X"02B4",
		X"0250",X"020A",X"019D",X"0152",X"00D6",X"0094",X"0043",X"FFF3",X"FF85",X"FF05",X"FEB6",X"FE35",X"FDB0",X"FD41",X"FCF1",X"FCB4",
		X"FCA1",X"FC97",X"FC9D",X"FCAB",X"FCB5",X"FC8D",X"FC39",X"FBC1",X"FB1A",X"FA5F",X"F9BA",X"F92B",X"F8D8",X"F8B2",X"F899",X"F89B",
		X"F8EF",X"F95A",X"F9D3",X"FA6B",X"FADE",X"FB56",X"FB76",X"FBC5",X"FBF7",X"FC3C",X"FC54",X"FC70",X"FCC6",X"FD37",X"FDDD",X"FE75",
		X"FF3F",X"FFE8",X"0090",X"0124",X"019F",X"0206",X"0258",X"026C",X"028C",X"02C2",X"0309",X"0349",X"0384",X"03C9",X"03FC",X"0420",
		X"0430",X"041D",X"03F7",X"03BC",X"0390",X"038E",X"03AA",X"03D9",X"0429",X"0491",X"051D",X"05B4",X"0642",X"0694",X"06FC",X"0745",
		X"074D",X"074C",X"0715",X"06DA",X"067D",X"0644",X"05FE",X"059C",X"0529",X"04AD",X"0438",X"03AB",X"031D",X"028A",X"01CD",X"00EC",
		X"FFEE",X"FF1B",X"FE63",X"FD9B",X"FD05",X"FCBA",X"FC7A",X"FC47",X"FC35",X"FC30",X"FC14",X"FBEA",X"FBAB",X"FB8E",X"FB50",X"FB25",
		X"FB34",X"FB22",X"FB28",X"FB37",X"FB76",X"FBCF",X"FC0C",X"FC48",X"FC9E",X"FD05",X"FD5A",X"FDB4",X"FDB7",X"FDBE",X"FDEE",X"FDE3",
		X"FDCC",X"FD90",X"FD59",X"FD2B",X"FCF4",X"FCDD",X"FCDE",X"FCEF",X"FD12",X"FD30",X"FD59",X"FD80",X"FDAB",X"FDED",X"FDEE",X"FDF9",
		X"FDFE",X"FDF6",X"FDFC",X"FE11",X"FE25",X"FE45",X"FE82",X"FEBC",X"FF0B",X"FF31",X"FF40",X"FF2C",X"FEE7",X"FE5F",X"FDDE",X"FD5D",
		X"FCDF",X"FC4A",X"FBD8",X"FB85",X"FB60",X"FB88",X"FBD8",X"FC6D",X"FD0B",X"FDA6",X"FE4F",X"FEBF",X"FF4B",X"FFDC",X"0026",X"0053",
		X"006A",X"0091",X"00E3",X"0147",X"01D6",X"0265",X"02EE",X"03A9",X"0452",X"0516",X"05DA",X"065D",X"06A6",X"06D8",X"06ED",X"06EF",
		X"070E",X"0732",X"0779",X"07BE",X"07F4",X"085B",X"08BE",X"090A",X"0945",X"097B",X"0990",X"0996",X"097F",X"0968",X"0925",X"08B1",
		X"0867",X"07D8",X"075A",X"06F2",X"0683",X"0634",X"05E5",X"0593",X"0551",X"0514",X"04D0",X"0480",X"042A",X"03BB",X"0315",X"0257",
		X"017B",X"0077",X"FF61",X"FE1F",X"FCC4",X"FB90",X"FA83",X"F9BD",X"F918",X"F8AC",X"F87B",X"F85B",X"F886",X"F8D5",X"F8FF",X"F91E",
		X"F937",X"F953",X"F956",X"F945",X"F90C",X"F8F6",X"F8DE",X"F8DB",X"F8DB",X"F905",X"F944",X"F973",X"F9A3",X"F9D3",X"FA02",X"FA11",
		X"FA11",X"F9F6",X"FA0F",X"FA23",X"FA25",X"FA1B",X"FA2D",X"FA52",X"FA93",X"FAF8",X"FB69",X"FBCA",X"FC57",X"FCEF",X"FD64",X"FDF4",
		X"FE51",X"FE8B",X"FE8A",X"FE95",X"FEB0",X"FEA8",X"FEA6",X"FEAC",X"FE94",X"FEAC",X"FEFD",X"FF64",X"FFCE",X"0040",X"00B1",X"0139",
		X"01BB",X"020B",X"0235",X"0241",X"022A",X"020B",X"01C4",X"017B",X"012B",X"00D7",X"00B1",X"0093",X"00AC",X"00CD",X"00F9",X"0134",
		X"0180",X"01D3",X"023E",X"0290",X"02CB",X"0306",X"0343",X"037D",X"03B2",X"03F1",X"0432",X"045F",X"047B",X"0496",X"0484",X"0481",
		X"047E",X"048F",X"04AE",X"04B6",X"04D0",X"04F6",X"050A",X"051E",X"051E",X"051C",X"050B",X"04E5",X"04E4",X"04BE",X"049E",X"0445",
		X"040B",X"03DC",X"03A8",X"039E",X"036C",X"0329",X"02FB",X"0298",X"0242",X"01DC",X"016E",X"00DB",X"002B",X"FFAF",X"FF39",X"FEF3",
		X"FECF",X"FEC5",X"FECE",X"FEEB",X"FF40",X"FFB4",X"0019",X"0086",X"00C2",X"00E4",X"00DC",X"00B0",X"0091",X"004E",X"0002",X"FF9E",
		X"FF21",X"FEC6",X"FE67",X"FE1F",X"FDFA",X"FDAF",X"FD67",X"FD3E",X"FCED",X"FCB0",X"FC7F",X"FC4C",X"FC19",X"FBE7",X"FBD1",X"FBD0",
		X"FBDE",X"FBDB",X"FBEC",X"FC1B",X"FC0D",X"FBF9",X"FC00",X"FBF5",X"FBCE",X"FBB6",X"FB9F",X"FB96",X"FB81",X"FBBE",X"FBF1",X"FC37",
		X"FCAE",X"FD11",X"FD95",X"FE0A",X"FE6E",X"FEC5",X"FF19",X"FF59",X"FF77",X"FF6E",X"FF51",X"FF40",X"FF37",X"FF1B",X"FF04",X"FEFA",
		X"FEE5",X"FE97",X"FE51",X"FE32",X"FE29",X"FDFE",X"FDF6",X"FE0D",X"FE53",X"FEC0",X"FF32",X"FFCA",X"004D",X"00EC",X"016F",X"01BB",
		X"021A",X"022B",X"0236",X"020A",X"01C9",X"018A",X"0144",X"0118",X"00DA",X"00B8",X"00AF",X"00CD",X"00F6",X"0121",X"0159",X"01A0",
		X"01D9",X"01F6",X"021C",X"0225",X"0247",X"0238",X"0235",X"021F",X"0205",X"021A",X"020E",X"01FD",X"01DC",X"01B9",X"016D",X"0120",
		X"00D4",X"00AC",X"006D",X"004F",X"003C",X"0057",X"0096",X"00CF",X"011A",X"0189",X"0203",X"0252",X"0290",X"02E1",X"0342",X"0385",
		X"03C2",X"03F7",X"0430",X"0457",X"0469",X"0489",X"049A",X"048D",X"047E",X"045C",X"043E",X"0419",X"03D4",X"038D",X"033C",X"02E7",
		X"02B9",X"028A",X"0261",X"020D",X"01CC",X"01B6",X"017C",X"0129",X"00BE",X"0047",X"FFE6",X"FF78",X"FEF6",X"FE5A",X"FDC2",X"FD59",
		X"FCF7",X"FCBB",X"FC91",X"FCA8",X"FCB8",X"FCC4",X"FCBF",X"FC85",X"FC60",X"FC14",X"FBAF",X"FB5F",X"FAFB",X"FA70",X"F9FF",X"F9A8",
		X"F9B6",X"F9BC",X"F9D7",X"FA06",X"FA26",X"FA65",X"FAC3",X"FB00",X"FAE0",X"FA9E",X"FA45",X"FA07",X"F9DC",X"F9CD",X"F9EA",X"FA5A",
		X"FAFD",X"FBDE",X"FCCA",X"FDCD",X"FEB8",X"FF64",X"FFD3",X"0020",X"0023",X"FFED",X"FFC3",X"FF8F",X"FF60",X"FF59",X"FF69",X"FF9B",
		X"0007",X"00B7",X"015C",X"01D4",X"0238",X"0261",X"0260",X"0237",X"01DC",X"0168",X"00DF",X"0064",X"0021",X"000D",X"002A",X"0086",
		X"00FD",X"0176",X"01DC",X"021B",X"026F",X"02A5",X"02BE",X"02A0",X"0263",X"0246",X"0262",X"0284",X"02E2",X"036B",X"03FA",X"0467",
		X"04C0",X"053B",X"0579",X"0589",X"057E",X"054F",X"04F5",X"04B8",X"049A",X"0478",X"044F",X"0440",X"046F",X"04B3",X"0508",X"0558",
		X"05A1",X"05CC",X"05E1",X"05E8",X"05C9",X"058A",X"0506",X"04D9",X"04AE",X"048C",X"047E",X"0460",X"0468",X"0481",X"0490",X"046C",
		X"040A",X"0380",X"02FE",X"022D",X"0174",X"00A7",X"FFA9",X"FED9",X"FE0B",X"FD6F",X"FCCB",X"FC64",X"FC3D",X"FBFF",X"FBD5",X"FB90",
		X"FB70",X"FB50",X"FB06",X"FAC5",X"FA89",X"FA39",X"F9F9",X"F9BA",X"F99A",X"F946",X"F917",X"F8F8",X"F89D",X"F828",X"F79D",X"F70F",
		X"F693",X"F63A",X"F615",X"F606",X"F600",X"F636",X"F68E",X"F726",X"F7E5",X"F895",X"F949",X"F9D5",X"FA65",X"FB1A",X"FBBD",X"FC6E",
		X"FD0D",X"FDC8",X"FE6B",X"FF35",X"0012",X"00C0",X"0166",X"01D0",X"023E",X"0297",X"02BE",X"02BC",X"027A",X"0230",X"0208",X"01F2",
		X"01D2",X"01C7",X"01CE",X"01DC",X"0217",X"027E",X"02DF",X"0311",X"0324",X"030D",X"02D8",X"0294",X"0259",X"0203",X"018B",X"0100",
		X"0086",X"0042",X"0016",X"000C",X"001E",X"0035",X"007F",X"00E3",X"0155",X"01C6",X"0226",X"0294",X"02DF",X"0302",X"0323",X"0337",
		X"0349",X"0365",X"0381",X"03AA",X"03C3",X"0409",X"0490",X"0535",X"05BA",X"0610",X"0654",X"0675",X"06A3",X"06BD",X"06AD",X"0671",
		X"062F",X"05E4",X"05A8",X"056D",X"0555",X"054D",X"0533",X"0534",X"051E",X"0537",X"0545",X"0552",X"0549",X"0527",X"04E8",X"04B0",
		X"046D",X"041E",X"03AB",X"0330",X"02BA",X"025A",X"01FE",X"018C",X"0143",X"0107",X"00F3",X"00B8",X"0047",X"FFDB",X"FF89",X"FF15",
		X"FE7B",X"FDB5",X"FCD8",X"FBE4",X"FAFD",X"FA14",X"F92B",X"F864",X"F7A9",X"F70B",X"F678",X"F643",X"F623",X"F604",X"F5CB",X"F590",
		X"F55C",X"F526",X"F4F9",X"F4B3",X"F489",X"F482",X"F48A",X"F4B9",X"F527",X"F5CE",X"F680",X"F749",X"F81C",X"F8C3",X"F97C",X"FA1C",
		X"FAA6",X"FB07",X"FB31",X"FB58",X"FB5E",X"FB49",X"FB8E",X"FBDB",X"FC6B",X"FCF1",X"FD6B",X"FE11",X"FEAD",X"FF7F",X"0047",X"00CB",
		X"0104",X"00F8",X"00DC",X"00AF",X"006B",X"0025",X"FFF3",X"FFF3",X"0026",X"0089",X"0141",X"0231",X"0328",X"0402",X"04A1",X"0518",
		X"0562",X"05A4",X"059E",X"058F",X"0571",X"0538",X"04E6",X"04DD",X"0517",X"056C",X"0602",X"0684",X"0707",X"0799",X"083C",X"08CB",
		X"091F",X"095A",X"0958",X"0955",X"0953",X"0982",X"0993",X"09A0",X"09D9",X"09EA",X"0A33",X"0A66",X"0A8F",X"0A7D",X"0A6D",X"0A1B",
		X"098B",X"08DC",X"0811",X"0770",X"06D3",X"062F",X"059D",X"0511",X"04BE",X"04A9",X"047A",X"046C",X"0464",X"0443",X"0429",X"041F",
		X"03F1",X"0383",X"02E8",X"024A",X"0190",X"00AB",X"FFC4",X"FEEA",X"FE2B",X"FD95",X"FD1E",X"FCB4",X"FC53",X"FC00",X"FBDA",X"FBB3",
		X"FB5E",X"FAF0",X"FA5A",X"F989",X"F88F",X"F78A",X"F694",X"F5AA",X"F4CC",X"F3D4",X"F31D",X"F2C3",X"F298",X"F2AC",X"F2DD",X"F345",
		X"F3C7",X"F453",X"F4F4",X"F582",X"F5DF",X"F633",X"F66D",X"F693",X"F6B9",X"F6DA",X"F715",X"F737",X"F770",X"F7A0",X"F7AC",X"F7A2",
		X"F76F",X"F760",X"F713",X"F6C1",X"F666",X"F5FA",X"F5E3",X"F5C2",X"F5D6",X"F61C",X"F685",X"F731",X"F817",X"F915",X"FA1B",X"FB3C",
		X"FC48",X"FD42",X"FE38",X"FF38",X"FFFB",X"00AB",X"0149",X"01D4",X"0255",X"02DD",X"0352",X"03F2",X"04A8",X"0542",X"05D9",X"0641",
		X"06B7",X"071C",X"0769",X"079F",X"078E",X"0776",X"0762",X"072F",X"0713",X"0735",X"0760",X"07A4",X"0803",X"0868",X"08EF",X"096F",
		X"0A1C",X"0AB3",X"0B1C",X"0B89",X"0BB7",X"0BBF",X"0BCD",X"0BE9",X"0C07",X"0C13",X"0C53",X"0CBF",X"0D27",X"0DA6",X"0E14",X"0E81",
		X"0ED3",X"0EF9",X"0EEF",X"0E7D",X"0DF8",X"0D3A",X"0C77",X"0BA0",X"0AC1",X"09E5",X"08FF",X"0850",X"07C5",X"0739",X"06BE",X"0627",
		X"059F",X"051C",X"049E",X"042A",X"035D",X"0296",X"01C3",X"00FF",X"003C",X"FF50",X"FE6D",X"FDA6",X"FCE1",X"FC4B",X"FBD3",X"FB45",
		X"FAB3",X"FA42",X"F9B6",X"F93D",X"F87D",X"F78E",X"F682",X"F56F",X"F45C",X"F33F",X"F237",X"F152",X"F0AD",X"F035",X"EFFA",X"EFDE",
		X"EFF1",X"F040",X"F08C",X"F0CE",X"F11B",X"F137",X"F142",X"F12B",X"F114",X"F111",X"F118",X"F11D",X"F12D",X"F171",X"F20C",X"F2D6",
		X"F3D4",X"F4F3",X"F61E",X"F730",X"F883",X"F9DA",X"FAED",X"FBBA",X"FC4B",X"FCCF",X"FD2D",X"FD91",X"FDE1",X"FE17",X"FE3B",X"FE5E",
		X"FEC2",X"FF42",X"FFC5",X"0043",X"00D7",X"0172",X"01EC",X"0262",X"02E8",X"0376",X"040A",X"045E",X"04BB",X"0514",X"0579",X"061E",
		X"06A8",X"0737",X"07C4",X"0879",X"0928",X"09B6",X"0A26",X"0A66",X"0A9B",X"0AA7",X"0A99",X"0A7D",X"0A61",X"0A2A",X"09E2",X"0988",
		X"0969",X"095C",X"0947",X"0937",X"092C",X"0945",X"0952",X"0986",X"09B1",X"09AF",X"09DA",X"0A03",X"09F6",X"09CD",X"0987",X"0957",
		X"0906",X"08D4",X"08A8",X"0859",X"0800",X"07B2",X"0787",X"077C",X"074F",X"06F8",X"06B7",X"063C",X"05DA",X"0534",X"043E",X"0327",
		X"01C4",X"0078",X"FF2F",X"FDE6",X"FCB1",X"FB95",X"FAA2",X"FA0A",X"F981",X"F943",X"F906",X"F8D3",X"F8AE",X"F895",X"F885",X"F83A",
		X"F7ED",X"F7A8",X"F762",X"F736",X"F707",X"F6C1",X"F6AB",X"F6B2",X"F6E7",X"F731",X"F756",X"F798",X"F7B8",X"F7C1",X"F7E3",X"F7DA",
		X"F7A6",X"F772",X"F744",X"F6FF",X"F6D9",X"F6B0",X"F690",X"F6BE",X"F6EB",X"F737",X"F7A4",X"F800",X"F86C",X"F8C7",X"F92F",X"F98E",
		X"F9FB",X"FA2D",X"FA5A",X"FA90",X"FAB6",X"FAC2",X"FA9F",X"FA98",X"FA9C",X"FA9F",X"FACB",X"FB27",X"FB8C",X"FC02",X"FC60",X"FCC1",
		X"FD01",X"FD2C",X"FD55",X"FD7A",X"FD53",X"FD1C",X"FCF9",X"FCE2",X"FCDD",X"FCDF",X"FD05",X"FD63",X"FDFA",X"FED4",X"FFC9",X"00CB",
		X"0207",X"0351",X"04AC",X"05D8",X"06DD",X"07CF",X"0896",X"094C",X"09ED",X"0A7F",X"0B15",X"0B8D",X"0C40",X"0D02",X"0DD4",X"0EA4",
		X"0F40",X"0FEE",X"106A",X"10C7",X"111D",X"111F",X"1102",X"10C4",X"1080",X"1035",X"0FCC",X"0F47",X"0EB7",X"0E3C",X"0DAF",X"0D2E",
		X"0CB0",X"0C2F",X"0B99",X"0ADF",X"0A54",X"09B3",X"0912",X"0838",X"074E",X"0670",X"0591",X"04B6",X"03DE",X"0305",X"022F",X"017E",
		X"00E6",X"004D",X"FF94",X"FEE5",X"FE1A",X"FD4D",X"FC92",X"FBD8",X"FB0A",X"FA50",X"F99B",X"F8ED",X"F86C",X"F7EE",X"F791",X"F766",
		X"F75E",X"F760",X"F760",X"F77C",X"F794",X"F7A9",X"F7A8",X"F77A",X"F734",X"F6E2",X"F680",X"F620",X"F5B3",X"F537",X"F4C4",X"F48C",
		X"F458",X"F449",X"F44B",X"F472",X"F4A0",X"F4E5",X"F511",X"F566",X"F5A0",X"F5D3",X"F618",X"F674",X"F6C1",X"F70E",X"F75E",X"F7A7",
		X"F7BE",X"F7EE",X"F81B",X"F847",X"F85A",X"F874",X"F8CB",X"F93D",X"F9A8",X"FA16",X"FA8C",X"FB07",X"FB6E",X"FBCA",X"FC34",X"FC85",
		X"FD11",X"FD95",X"FE26",X"FEAB",X"FF3C",X"FFC7",X"007B",X"011F",X"01A7",X"020D",X"027F",X"02DA",X"031D",X"0383",X"03C7",X"040E",
		X"044E",X"04B1",X"053A",X"059C",X"0621",X"068D",X"06F4",X"0742",X"0791",X"079C",X"0788",X"0775",X"0747",X"071F",X"0704",X"0709",
		X"0703",X"0707",X"0727",X"0771",X"07A7",X"07BF",X"07E2",X"07F5",X"07F3",X"07EE",X"07E4",X"07B5",X"076E",X"0733",X"072B",X"0704",
		X"06D5",X"06A5",X"0668",X"0646",X"05FB",X"05AE",X"051E",X"048F",X"03F1",X"0361",X"02F3",X"0284",X"022C",X"0220",X"0263",X"02AA",
		X"031C",X"0380",X"0413",X"04A7",X"052D",X"057B",X"05BF",X"05D8",X"05B5",X"0583",X"052B",X"04B4",X"040F",X"037E",X"02A7",X"01D7",
		X"0100",X"0009",X"FF22",X"FE36",X"FD73",X"FCD5",X"FC6E",X"FC1B",X"FBEF",X"FBBC",X"FBC2",X"FBC3",X"FBEA",X"FBF6",X"FBD9",X"FB9E",
		X"FB51",X"FB05",X"FAA4",X"FA5A",X"FA04",X"F9DE",X"F99B",X"F9A8",X"F9B2",X"F9F2",X"FA0A",X"FA15",X"FA26",X"FA2C",X"FA2E",X"FA10",
		X"F9E7",X"F991",X"F947",X"F90C",X"F8F3",X"F8DB",X"F8E2",X"F910",X"F957",X"F9B3",X"FA08",X"FA56",X"FA97",X"FAF9",X"FB48",X"FB72",
		X"FB8F",X"FB51",X"FAF8",X"FAB7",X"FA9D",X"FA76",X"FA45",X"FA20",X"FA20",X"FA50",X"FAAF",X"FB25",X"FB91",X"FBF4",X"FC64",X"FCA8",
		X"FCF3",X"FD3A",X"FD65",X"FD71",X"FD77",X"FDAD",X"FE02",X"FE62",X"FEB7",X"FF33",X"FFD1",X"0072",X"011E",X"01CA",X"0286",X"0321",
		X"03AE",X"0432",X"0483",X"04D3",X"04EE",X"0527",X"052A",X"051A",X"04F9",X"04A6",X"0495",X"048D",X"0468",X"0418",X"03D0",X"03A4",
		X"037F",X"0369",X"0365",X"0343",X"033C",X"0368",X"03AC",X"0407",X"047A",X"0524",X"059C",X"05CE",X"062F",X"068A",X"06F0",X"071D",
		X"0734",X"071E",X"06E4",X"069D",X"063B",X"05D6",X"0560",X"04D2",X"044C",X"03E6",X"03AB",X"03AC",X"03B8",X"03E8",X"0444",X"04A7",
		X"0519",X"058A",X"05E1",X"063E",X"069C",X"06FD",X"0739",X"0767",X"0797",X"079B",X"07A5",X"07B3",X"07B1",X"07C0",X"07BA",X"079E",
		X"0764",X"0710",X"0692",X"0606",X"056C",X"04CC",X"03F9",X"033B",X"024A",X"0168",X"009E",X"FFF4",X"FF3A",X"FE5E",X"FD86",X"FCB3",
		X"FBEB",X"FB26",X"FA75",X"F9C1",X"F908",X"F824",X"F72B",X"F677",X"F5E9",X"F55C",X"F4EE",X"F45B",X"F3DC",X"F373",X"F2F5",X"F27A",
		X"F1EC",X"F154",X"F09E",X"EFDD",X"EF52",X"EEEC",X"EEA5",X"EE9A",X"EED2",X"EF2E",X"EFCB",X"F08B",X"F18E",X"F27E",X"F353",X"F422",
		X"F4DE",X"F561",X"F5CA",X"F629",X"F687",X"F6CE",X"F70A",X"F76F",X"F7DE",X"F886",X"F931",X"F9BC",X"FA1D",X"FA7B",X"FAD7",X"FB30",
		X"FB7C",X"FBBB",X"FBE0",X"FBE0",X"FBD3",X"FC12",X"FC99",X"FD45",X"FE19",X"FEFF",X"0013",X"0162",X"02F5",X"0459",X"0585",X"068A",
		X"0770",X"082C",X"08E7",X"0992",X"0A05",X"0A73",X"0ABF",X"0B0E",X"0B9B",X"0C44",X"0CF5",X"0D8C",X"0E2C",X"0EE1",X"0F8B",X"1036",
		X"10DB",X"112D",X"1167",X"1168",X"113D",X"10F2",X"10A2",X"106B",X"1022",X"0FEE",X"0FE7",X"0FE7",X"101B",X"1068",X"10D1",X"114F",
		X"1172",X"11A5",X"11B9",X"11BF",X"117C",X"1114",X"10A2",X"1007",X"0F72",X"0EC0",X"0E19",X"0D73",X"0CC9",X"0BEF",X"0AFC",X"09FC",
		X"08EB",X"0790",X"061B",X"04A2",X"030D",X"0195",X"0021",X"FED5",X"FD8F",X"FC8F",X"FBD0",X"FB62",X"FB1A",X"FAD4",X"FAAA",X"FA85",
		X"FA5B",X"FA21",X"F9B5",X"F931",X"F87F",X"F7AD",X"F6B7",X"F596",X"F468",X"F34B",X"F257",X"F181",X"F0DD",X"F052",X"EFF3",X"EFD2",
		X"EFED",X"F00E",X"F002",X"EFEE",X"EFC5",X"EF69",X"EF0D",X"EEB8",X"EE71",X"EE00",X"ED9D",X"ED63",X"ED5F",X"ED5E",X"ED79",X"EDC8",
		X"EE02",X"EE6F",X"EEED",X"EF8C",X"F027",X"F0F1",X"F199",X"F232",X"F291",X"F306",X"F387",X"F400",X"F48F",X"F508",X"F5A1",X"F641",
		X"F6D6",X"F79D",X"F865",X"F8F7",X"F957",X"F9A5",X"F9E5",X"FA1A",X"FA3E",X"FA55",X"FA66",X"FAA2",X"FB1C",X"FB98",X"FC4D",X"FD0D",
		X"FE03",X"FF2C",X"0048",X"016E",X"0286",X"03A4",X"04D3",X"05C0",X"066E",X"06F0",X"0759",X"07A2",X"07EF",X"0833",X"0890",X"08ED",
		X"0967",X"09DF",X"0A75",X"0AF3",X"0B98",X"0C20",X"0CB0",X"0D29",X"0D7D",X"0DB6",X"0DB0",X"0DC3",X"0DDD",X"0E09",X"0E28",X"0E19",
		X"0DDD",X"0DCA",X"0DDE",X"0E07",X"0E0C",X"0E16",X"0E31",X"0E33",X"0E44",X"0E4C",X"0E51",X"0E88",X"0EA5",X"0ED0",X"0EF4",X"0F3F",
		X"0F7E",X"0FBC",X"0FFA",X"1022",X"1015",X"0FE5",X"0F80",X"0F17",X"0E97",X"0DF1",X"0D1D",X"0C0C",X"0AF9",X"09C8",X"089E",X"0753",
		X"0604",X"04CC",X"0395",X"0283",X"01AA",X"00C1",X"0025",X"FFC1",X"FF5B",X"FF07",X"FE9E",X"FE2C",X"FDAD",X"FD20",X"FC74",X"FBA9",
		X"FAD3",X"F9F0",X"F930",X"F874",X"F7CB",X"F71A",X"F675",X"F5E9",X"F5A5",X"F576",X"F552",X"F531",X"F4F8",X"F4C7",X"F49E",X"F465",
		X"F414",X"F3BB",X"F363",X"F31F",X"F2D5",X"F29D",X"F296",X"F2B4",X"F2C9",X"F317",X"F357",X"F386",X"F3AE",X"F3B9",X"F3DF",X"F3F0",
		X"F404",X"F3F3",X"F3AD",X"F38E",X"F384",X"F3A8",X"F3C8",X"F3ED",X"F40D",X"F47F",X"F523",X"F5C2",X"F644",X"F6B8",X"F702",X"F74A",
		X"F781",X"F794",X"F7A1",X"F79C",X"F7AB",X"F7AC",X"F7F1",X"F869",X"F8FA",X"F992",X"FA53",X"FB3A",X"FC1D",X"FCE9",X"FD8E",X"FE22",
		X"FEAA",X"FF16",X"FF50",X"FF73",X"FFA1",X"FFFC",X"006B",X"010E",X"01D8",X"0295",X"0380",X"048B",X"05B3",X"06DC",X"07D8",X"08AB",
		X"0966",X"09FD",X"0A84",X"0AF5",X"0B42",X"0B87",X"0BBA",X"0BEF",X"0C25",X"0C7C",X"0CE1",X"0D41",X"0DAF",X"0DFE",X"0E43",X"0E7D",
		X"0EB5",X"0EF8",X"0F39",X"0F3C",X"0F1A",X"0EE5",X"0EA3",X"0E66",X"0E3F",X"0E15",X"0DDB",X"0DA0",X"0D88",X"0D93",X"0DC4",X"0DDC",
		X"0DC8",X"0D8B",X"0D57",X"0D01",X"0C99",X"0C0F",X"0B66",X"0ACC",X"0A19",X"0977",X"08E5",X"0848",X"07A0",X"0707",X"065E",X"05AF",
		X"04D3",X"03F7",X"0313",X"0212",X"0114",X"0014",X"FF1C",X"FE55",X"FD8E",X"FCD4",X"FC1D",X"FB4C",X"FA91",X"F9B2",X"F8D3",X"F7DD",
		X"F6E0",X"F60F",X"F540",X"F48F",X"F40B",X"F39B",X"F338",X"F2F1",X"F2AE",X"F271",X"F22D",X"F1F8",X"F19D",X"F13E",X"F10F",X"F0BD",
		X"F08E",X"F047",X"F030",X"F035",X"F04A",X"F076",X"F09B",X"F0C7",X"F0EB",X"F106",X"F0FB",X"F0DF",X"F09C",X"F05C",X"F029",X"F003",
		X"F016",X"F04F",X"F0AB",X"F15F",X"F238",X"F32E",X"F433",X"F534",X"F640",X"F72D",X"F7F1",X"F889",X"F915",X"F992",X"FA11",X"FAB7",
		X"FB5D",X"FBFB",X"FCA8",X"FD7F",X"FE5D",X"FF81",X"009A",X"018D",X"029A",X"036D",X"0467",X"0544",X"05D5",X"066A",X"06D7",X"070B",
		X"0733",X"0753",X"0764",X"0791",X"07D8",X"083D",X"088F",X"090A",X"096D",X"09B2",X"09F0",X"0A02",X"09F1",X"09CC",X"099E",X"0992",
		X"099D",X"09D7",X"0A15",X"0A47",X"0AA6",X"0AFF",X"0B89",X"0BDD",X"0C0A",X"0C22",X"0C15",X"0BEB",X"0BAF",X"0B70",X"0B13",X"0AD6",
		X"0AA2",X"0A93",X"0A88",X"0A70",X"0A6B",X"0A79",X"0A9D",X"0A90",X"0A99",X"0A9A",X"0A66",X"0A0A",X"099E",X"0913",X"0880",X"07EB",
		X"0736",X"067D",X"05F4",X"0578",X"04F6",X"0484",X"0432",X"03D5",X"0387",X"0344",X"02F6",X"02E1",X"02AD",X"025B",X"01D8",X"014B",
		X"009D",X"FFF5",X"FF3E",X"FE86",X"FDD3",X"FD47",X"FCC8",X"FC57",X"FC41",X"FBE6",X"FB93",X"FB34",X"FAD4",X"FA63",X"F9C9",X"F91B",
		X"F868",X"F7E2",X"F76D",X"F705",X"F68F",X"F649",X"F609",X"F5D1",X"F5C5",X"F599",X"F552",X"F52A",X"F52B",X"F50F",X"F507",X"F4D8",
		X"F4BA",X"F49E",X"F4AB",X"F4C9",X"F4DC",X"F4FD",X"F50D",X"F549",X"F5AB",X"F627",X"F68D",X"F6D1",X"F714",X"F76A",X"F7B6",X"F809",
		X"F855",X"F8B0",X"F934",X"F9B0",X"FA3C",X"FAEF",X"FB66",X"FBE8",X"FC54",X"FCB2",X"FD0A",X"FD3C",X"FD6D",X"FD8C",X"FDB6",X"FDE7",
		X"FDF6",X"FDE8",X"FDDF",X"FDB7",X"FD9F",X"FD9D",X"FDA6",X"FDEC",X"FE3A",X"FE77",X"FF00",X"FFBB",X"005B",X"00E4",X"0177",X"021F",
		X"02A0",X"0319",X"0392",X"0400",X"0478",X"04E7",X"0550",X"05AC",X"0611",X"0648",X"0681",X"06A9",X"06AD",X"06BD",X"06E0",X"0709",
		X"073D",X"077E",X"07D8",X"084D",X"08D3",X"0978",X"09EE",X"0A4F",X"0AA0",X"0ACF",X"0AE3",X"0AF5",X"0AD9",X"0AAB",X"0A84",X"0A5B",
		X"0A40",X"0A18",X"09E4",X"09DE",X"09D3",X"09DC",X"09DB",X"09C4",X"0990",X"095B",X"0910",X"08D5",X"086A",X"07EB",X"0788",X"0727",
		X"06DB",X"0684",X"0634",X"05E4",X"05A7",X"054F",X"050D",X"04A0",X"0437",X"03C5",X"0355",X"02D7",X"022F",X"0185",X"00A5",X"FFC1",
		X"FEE4",X"FE00",X"FD31",X"FC6A",X"FBBE",X"FB28",X"FAA8",X"FA4D",X"F9F1",X"F9AA",X"F96C",X"F92F",X"F8FC",X"F901",X"F8E5",X"F8CB",
		X"F8B4",X"F8AA",X"F8A8",X"F89D",X"F8A1",X"F86E",X"F862",X"F854",X"F818",X"F7C7",X"F773",X"F721",X"F6E0",X"F6C0",X"F6C0",X"F6B0",
		X"F694",X"F6AB",X"F6C2",X"F6F3",X"F704",X"F6E4",X"F6D9",X"F6D7",X"F6D7",X"F6A7",X"F696",X"F692",X"F697",X"F6EB",X"F74C",X"F7C5",
		X"F82C",X"F8C3",X"F980",X"FA38",X"FAB0",X"FAFE",X"FB2F",X"FB28",X"FAF8",X"FA9D",X"FA40",X"FA12",X"FA21",X"FA45",X"FAA5",X"FB1D",
		X"FBA2",X"FC4C",X"FCD0",X"FD4C",X"FD9B",X"FDAF",X"FDF9",X"FE12",X"FE57",X"FEAC",X"FF32",X"FFF8",X"00CD",X"01CB",X"02E8",X"03E1",
		X"04F2",X"060D",X"06DF",X"0773",X"07D1",X"0813",X"0842",X"0864",X"0874",X"087A",X"0884",X"0898",X"08A1",X"0910",X"09A7",X"0A28",
		X"0A89",X"0AC5",X"0B01",X"0B68",X"0BB7",X"0BE4",X"0BD8",X"0BB3",X"0BA5",X"0B9C",X"0BC1",X"0BE6",X"0BF8",X"0BDE",X"0BCC",X"0BA0",
		X"0B64",X"0B0D",X"0A99",X"09F1",X"0939",X"08A2",X"081F",X"0779",X"06DA",X"0642",X"058E",X"04DE",X"0440",X"03B8",X"0323",X"02A7",
		X"0239",X"01D6",X"01A1",X"0144",X"0121",X"00FF",X"00D8",X"00B7",X"0064",X"FFF5",X"FFAF",X"FF5E",X"FF0E",X"FEA6",X"FE28",X"FDB1",
		X"FD35",X"FCF1",X"FCB1",X"FC89",X"FC30",X"FBD9",X"FBA2",X"FB68",X"FB0D",X"FAB0",X"FA28",X"F98B",X"F8EC",X"F851",X"F7A9",X"F6FD",
		X"F66F",X"F5EC",X"F55E",X"F4E6",X"F48E",X"F446",X"F3F8",X"F3AC",X"F337",X"F2E0",X"F27F",X"F268",X"F264",X"F256",X"F2A2",X"F2D9",
		X"F338",X"F3AA",X"F41A",X"F48B",X"F52D",X"F5B5",X"F63C",X"F6B6",X"F720",X"F779",X"F7AA",X"F7CE",X"F7E2",X"F803",X"F84C",X"F8B7",
		X"F943",X"F9D0",X"FA82",X"FB4E",X"FC49",X"FD34",X"FE4F",X"FF45",X"0024",X"0108",X"01D4",X"0295",X"0359",X"040E",X"04D3",X"05C1",
		X"0682",X"0757",X"081B",X"08E4",X"098F",X"0A3B",X"0AAE",X"0AEF",X"0B17",X"0B1C",X"0B08",X"0AD5",X"0A85",X"0A20",X"09B6",X"0982",
		X"0963",X"0949",X"0954",X"0948",X"095F",X"096C",X"098D",X"09A1",X"09C3",X"0995",X"096C",X"091E",X"08C7",X"0893",X"082E",X"07CC",
		X"0748",X"06CB",X"064B",X"05DD",X"0570",X"0501",X"0472",X"040C",X"0389",X"032F",X"02EF",X"02C1",X"02AD",X"0298",X"02AA",X"02CC",
		X"02EC",X"02FC",X"030F",X"031C",X"030D",X"02EF",X"02B7",X"0242",X"01B8",X"0130",X"00CC",X"0060",X"FFFD",X"FF9D",X"FF71",X"FF67",
		X"FF3C",X"FEF5",X"FEB8",X"FE93",X"FE6A",X"FE34",X"FDEE",X"FD98",X"FD1D",X"FCB7",X"FC3A",X"FBD6",X"FB7A",X"FB2A",X"FAFB",X"FAB8",
		X"FA9E",X"FAB5",X"FAEC",X"FB1D",X"FB30",X"FB37",X"FB3D",X"FB2E",X"FB12",X"FACA",X"FA5E",X"FA23",X"F9CE",X"F982",X"F94E",X"F90C",
		X"F8CD",X"F899",X"F868",X"F83D",X"F82D",X"F813",X"F827",X"F834",X"F849",X"F85E",X"F88C",X"F8DB",X"F91E",X"F97A",X"F9D5",X"FA33",
		X"FA7F",X"FB10",X"FB93",X"FBF1",X"FC2E",X"FC5D",X"FC8E",X"FCC5",X"FCEE",X"FCFF",X"FD08",X"FCFA",X"FD16",X"FD40",X"FD58",X"FD88",
		X"FDA2",X"FDD8",X"FE0B",X"FE3D",X"FE7A",X"FEAC",X"FEF1",X"FF6F",X"FFFB",X"0089",X"00FF",X"0150",X"01A1",X"01A9",X"0191",X"0149",
		X"00FF",X"00B0",X"009F",X"00D1",X"00F8",X"016C",X"0229",X"02E1",X"03D3",X"048B",X"052D",X"0590",X"0593",X"0591",X"055A",X"04FF",
		X"0497",X"0451",X"0443",X"046D",X"04B5",X"053E",X"05C9",X"069A",X"0793",X"0889",X"0981",X"09EF",X"0A42",X"0A8D",X"0AB6",X"0AB2",
		X"0A86",X"0A45",X"09E9",X"09B2",X"0997",X"09A8",X"09B9",X"09C9",X"09CC",X"09B3",X"09BB",X"0990",X"0951",X"0902",X"08B4",X"083D",
		X"0808",X"07DB",X"07CE",X"07AC",X"0758",X"072C",X"06FA",X"0697",X"0607",X"0546",X"0476",X"03A6",X"029F",X"019E",X"008C",X"FF75",
		X"FE7F",X"FDCB",X"FD18",X"FC64",X"FBBF",X"FB35",X"FAF1",X"FA90",X"FA1D",X"F998",X"F8F4",X"F869",X"F7C3",X"F71A",X"F680",X"F5F1",
		X"F586",X"F51D",X"F4BA",X"F489",X"F45E",X"F42B",X"F3F2",X"F3B6",X"F374",X"F35F",X"F34E",X"F366",X"F34D",X"F33F",X"F333",X"F2FD",
		X"F2B4",X"F2A1",X"F285",X"F22F",X"F1E7",X"F1A0",X"F19E",X"F1A5",X"F1D8",X"F23E",X"F2AD",X"F33D",X"F3FC",X"F4D6",X"F5AE",X"F699",
		X"F768",X"F835",X"F8F9",X"F9C4",X"FA56",X"FAE2",X"FB47",X"FBAB",X"FC1E",X"FC68",X"FCD0",X"FD17",X"FD69",X"FDD6",X"FE59",X"FEFE",
		X"FF84",X"0019",X"00E3",X"0184",X"024F",X"0335",X"042B",X"052C",X"061D",X"06EE",X"07CF",X"0893",X"0962",X"0A17",X"0AA6",X"0B29",
		X"0BAE",X"0C44",X"0CCB",X"0D46",X"0DC5",X"0E2D",X"0E73",X"0EC6",X"0F16",X"0F5C",X"0F89",X"0F7B",X"0F64",X"0F49",X"0F09",X"0EA4",
		X"0E0E",X"0D54",X"0C7F",X"0BBD",X"0B14",X"0A97",X"0A41",X"0A08",X"09D0",X"09C1",X"09C0",X"09CA",X"09B8",X"09A0",X"096A",X"0932",
		X"0914",X"08DE",X"08B6",X"0888",X"0877",X"0855",X"080D",X"07C6",X"0783",X"0734",X"06D1",X"061A",X"055A",X"049C",X"03C1",X"02DE",
		X"01F0",X"00CF",X"FFEC",X"FF3B",X"FEBA",X"FE53",X"FDFB",X"FDDB",X"FDD5",X"FE00",X"FE11",X"FDF0",X"FDA0",X"FD35",X"FCC3",X"FC3C",
		X"FBBD",X"FB4A",X"FAB8",X"FA72",X"FA41",X"FA29",X"F9FE",X"F9BB",X"F98B",X"F93A",X"F8B3",X"F7EA",X"F714",X"F627",X"F52D",X"F476",
		X"F3A8",X"F2BF",X"F1F0",X"F112",X"F079",X"F005",X"EFA8",X"EF53",X"EEFF",X"EEA8",X"EE4C",X"EE04",X"EDAA",X"ED41",X"ECD6",X"EC6D",
		X"EC1A",X"EC0C",X"EC19",X"EC6A",X"ECF0",X"EDB8",X"EEAA",X"EFB7",X"F0E0",X"F1F8",X"F2F1",X"F3E2",X"F4C1",X"F597",X"F66A",X"F734",
		X"F814",X"F902",X"F9E9",X"FAC5",X"FBB9",X"FCDD",X"FE20",X"FF6F",X"00BF",X"01F8",X"0337",X"04A6",X"060D",X"0735",X"0833",X"08EC",
		X"096D",X"09FD",X"0A86",X"0ADE",X"0B1C",X"0B7E",X"0C01",X"0C73",X"0D07",X"0D9E",X"0E30",X"0EC2",X"0F6D",X"100B",X"108E",X"1107",
		X"115E",X"11B0",X"1203",X"1240",X"122B",X"11F8",X"11C3",X"117E",X"1121",X"10AF",X"101B",X"0F92",X"0F16",X"0E95",X"0DF2",X"0D29",
		X"0C6F",X"0BBA",X"0B04",X"0A4D",X"09A8",X"08FA",X"0832",X"07A1",X"0728",X"06D8",X"069B",X"0657",X"0616",X"05C0",X"0591",X"0563",
		X"0513",X"048F",X"040C",X"038F",X"02F4",X"026A",X"01F1",X"016F",X"0119",X"00E3",X"00CA",X"00B1",X"00A2",X"0097",X"0090",X"0065",
		X"0005",X"FF45",X"FE4C",X"FD20",X"FBC3",X"FA64",X"F900",X"F7B5",X"F6A2",X"F5C9",X"F541",X"F4F8",X"F4EC",X"F532",X"F577",X"F5E3",
		X"F639",X"F684",X"F6C3",X"F6E0",X"F70B",X"F759",X"F794",X"F7BA",X"F7E8",X"F80E",X"F84B",X"F886",X"F8ED",X"F967",X"F9A6",X"F9E0",
		X"FA2C",X"FA56",X"FA75",X"FA91",X"FA76",X"FA35",X"F9EF",X"F97C",X"F8F4",X"F875",X"F811",X"F7D1",X"F767",X"F715",X"F6E4",X"F6C7",
		X"F6D5",X"F6E4",X"F6E9",X"F719",X"F787",X"F7F1",X"F846",X"F89E",X"F8FA",X"F955",X"F988",X"F9A0",X"F9E3",X"FA12",X"FA66",X"FAD2",
		X"FB1D",X"FB86",X"FBCE",X"FC2E",X"FC86",X"FCDD",X"FD3B",X"FD80",X"FDB6",X"FDFB",X"FE3F",X"FE7B",X"FEBF",X"FF1E",X"FF83",X"FFCD",
		X"0034",X"006F",X"00D5",X"012B",X"016E",X"01C6",X"0228",X"028B",X"02F3",X"0383",X"0422",X"04B8",X"0549",X"05EE",X"0687",X"0730",
		X"07D8",X"08AD",X"0965",X"0A29",X"0AE3",X"0B93",X"0C2D",X"0CB6",X"0CFE",X"0D3C",X"0D51",X"0D2D",X"0D0C",X"0CCA",X"0C82",X"0C47",
		X"0BFE",X"0BBF",X"0B8B",X"0B46",X"0B1E",X"0AD9",X"0A8D",X"0A5F",X"0A11",X"098F",X"08E3",X"0806",X"0718",X"05FD",X"04E3",X"03BF",
		X"02A4",X"019A",X"00C5",X"0030",X"FFA5",X"FF3F",X"FEFC",X"FEB6",X"FE94",X"FE6C",X"FE66",X"FE62",X"FE5B",X"FE6D",X"FE49",X"FE32",
		X"FDF2",X"FDCC",X"FDBF",X"FD87",X"FD40",X"FCF5",X"FC9A",X"FC2A",X"FBD9",X"FB7D",X"FB03",X"FA83",X"FA0B",X"F9CC",X"F984",X"F94C",
		X"F927",X"F937",X"F97E",X"F9D2",X"FA3C",X"FAC7",X"FB4B",X"FBA5",X"FBFB",X"FC31",X"FC59",X"FC85",X"FC9B",X"FCAC",X"FCD4",X"FD04",
		X"FD35",X"FD78",X"FDB9",X"FE16",X"FE86",X"FEBD",X"FF0F",X"FF5D",X"FFA0",X"FFB0",X"FFBF",X"FFB3",X"FF73",X"FF29",X"FEE8",X"FEA5",
		X"FE44",X"FDFD",X"FDCE",X"FDB7",X"FDF6",X"FE4D",X"FE90",X"FEBA",X"FED5",X"FED7",X"FEE8",X"FED9",X"FEC4",X"FE6F",X"FE12",X"FDBF",
		X"FD4F",X"FD1C",X"FCE0",X"FCB8",X"FC93",X"FC99",X"FCB2",X"FCE8",X"FD3D",X"FD95",X"FDD9",X"FE3D",X"FE68",X"FE8A",X"FEB5",X"FEC2",
		X"FEED",X"FF1B",X"FF40",X"FF4E",X"FF59",X"FF89",X"FFC9",X"FFE2",X"FFFA",X"FFFD",X"0007",X"0005",X"002A",X"0046",X"0064",X"008D",
		X"00C7",X"011A",X"017B",X"01F5",X"027D",X"02F3",X"0332",X"038F",X"03F5",X"0448",X"049E",X"04EF",X"053B",X"0582",X"05B1",X"05EA",
		X"062F",X"0660",X"0688",X"06B7",X"06E6",X"0708",X"0729",X"0755",X"077B",X"079A",X"0774",X"0743",X"06EB",X"0689",X"0616",X"058E",
		X"04E3",X"043C",X"03A4",X"02FD",X"0260",X"01B8",X"0101",X"0052",X"FFD4",X"FF7C",X"FF37",X"FF18",X"FF2B",X"FF51",X"FF8B",X"FFC8",
		X"FFFE",X"0021",X"0003",X"FFD0",X"FF7F",X"FF2F",X"FEBE",X"FE38",X"FDC9",X"FD70",X"FD19",X"FCFD",X"FCE7",X"FCD0",X"FCD3",X"FCCE",
		X"FCF7",X"FD01",X"FD18",X"FD06",X"FCFA",X"FCC6",X"FC6B",X"FC18",X"FBCF",X"FB81",X"FB2F",X"FB1C",X"FB13",X"FB26",X"FB67",X"FBBF",
		X"FC31",X"FC9D",X"FCFB",X"FD5E",X"FDBC",X"FE14",X"FE30",X"FE73",X"FE8F",X"FE9C",X"FE91",X"FE73",X"FE61",X"FE40",X"FE4B",X"FE6D",
		X"FE78",X"FE77",X"FE7D",X"FE91",X"FEDB",X"FF38",X"FF75",X"FF91",X"FFBF",X"FFBE",X"FFB9",X"FF97",X"FF6B",X"FF27",X"FEE9",X"FEA1",
		X"FE5A",X"FE2D",X"FE14",X"FE03",X"FDF8",X"FE01",X"FDFE",X"FE1B",X"FE26",X"FE3D",X"FE3D",X"FE47",X"FE40",X"FE06",X"FDDC",X"FDA8",
		X"FD91",X"FDB0",X"FDEA",X"FE39",X"FE8B",X"FF02",X"FF95",X"001B",X"0086",X"00FB",X"0168",X"01B0",X"01B4",X"01AD",X"01A0",X"018A",
		X"0187",X"01A4",X"01D5",X"01F9",X"023F",X"0293",X"0300",X"0353",X"03A9",X"03EF",X"0428",X"045C",X"046C",X"045A",X"042C",X"03B7",
		X"0373",X"0341",X"031D",X"033A",X"0353",X"03A6",X"03E6",X"0444",X"0489",X"04C9",X"0513",X"0548",X"0568",X"056A",X"0577",X"0570",
		X"0561",X"0533",X"04F2",X"047E",X"0412",X"03B7",X"0349",X"02DA",X"0274",X"01FE",X"01A1",X"0144",X"00C8",X"0043",X"FF81",X"FEB4",
		X"FDC2",X"FCED",X"FC3B",X"FB7D",X"FAC6",X"FA49",X"FA05",X"F9F7",X"FA0D",X"FA06",X"FA33",X"FA41",X"FA4C",X"FA7A",X"FAAE",X"FAC6",
		X"FAC2",X"FAA7",X"FA9B",X"FA8E",X"FA89",X"FA97",X"FA7A",X"FA84",X"FABC",X"FAF1",X"FB51",X"FBA9",X"FC1A",X"FC9F",X"FD2F",X"FDC0",
		X"FE21",X"FE61",X"FE90",X"FEB4",X"FEE0",X"FF44",X"FF83",X"FFD6",X"002C",X"00C2",X"015B",X"020F",X"02CF",X"0379",X"0406",X"0481",
		X"0507",X"0565",X"05A5",X"05C8",X"05D7",X"05D8",X"05D2",X"05CB",X"05DC",X"05D5",X"05D6",X"05F1",X"0609",X"0603",X"05D6",X"05B5",
		X"0588",X"052A",X"04AD",X"0449",X"03BE",X"0331",X"02CE",X"0251",X"01DE",X"0176",X"0113",X"00D3",X"0080",X"0005",X"FF97",X"FEF6",
		X"FE67",X"FDBD",X"FD06",X"FC5F",X"FBBF",X"FB56",X"FB23",X"FB04",X"FB0F",X"FB5F",X"FBB3",X"FC2A",X"FC9C",X"FD16",X"FD8B",X"FDDC",
		X"FE20",X"FE59",X"FE82",X"FE94",X"FEA4",X"FEC6",X"FEF2",X"FF51",X"FF95",X"FFB5",X"FFD2",X"FFD9",X"FFBE",X"FF9A",X"FF5D",X"FF1E",
		X"FED7",X"FE8A",X"FE6A",X"FE5D",X"FE97",X"FED6",X"FF4D",X"FFBC",X"0022",X"00A0",X"010D",X"0140",X"0160",X"0170",X"016A",X"0170",
		X"015B",X"012E",X"00E6",X"00C2",X"00A2",X"0087",X"0067",X"006D",X"0060",X"0053",X"0023",X"FFEA",X"FFAE",X"FF38",X"FEB5",X"FE28",
		X"FDA8",X"FD2C",X"FCD7",X"FC8C",X"FC7A",X"FC97",X"FCD8",X"FD1D",X"FD83",X"FDEA",X"FE2B",X"FE6E",X"FEA4",X"FEC5",X"FEF2",X"FF1B",
		X"FF5C",X"FF9C",X"FFE0",X"004B",X"00A6",X"0117",X"018E",X"01D6",X"020F",X"023E",X"0249",X"021E",X"01B8",X"012D",X"0092",X"0013",
		X"FF89",X"FF38",X"FF2D",X"FF47",X"FF50",X"FF91",X"FFEE",X"0056",X"00E2",X"0148",X"01A0",X"01DE",X"021F",X"0249",X"0274",X"02A8",
		X"02C2",X"02BF",X"02B4",X"02A7",X"0279",X"021C",X"01BA",X"0143",X"00FC",X"00AE",X"0072",X"002F",X"FFFD",X"FFDB",X"FFB8",X"FF9F",
		X"FF9D",X"FF8B",X"FF5E",X"FF2F",X"FF11",X"FEFB",X"FEED",X"FEDF",X"FEFA",X"FF23",X"FF28",X"FF43",X"FF67",X"FF79",X"FF72",X"FF5D",
		X"FF1F",X"FED9",X"FE80",X"FE38",X"FDFC",X"FDCE",X"FDCA",X"FDDE",X"FDF1",X"FE2D",X"FE92",X"FF19",X"FFAF",X"0025",X"0046",X"003E",
		X"002E",X"FFE9",X"FF65",X"FEBE",X"FE2B",X"FD7D",X"FCDC",X"FC6D",X"FC03",X"FBD0",X"FBB9",X"FBC8",X"FBDE",X"FBFF",X"FC52",X"FCBD",
		X"FD27",X"FD9B",X"FDD7",X"FDF4",X"FE13",X"FE40",X"FE8C",X"FEBD",X"FEEE",X"FF3E",X"FFA9",X"002B",X"0097",X"00DF",X"010E",X"0112",
		X"00FA",X"00CB",X"0070",X"FFF2",X"FF98",X"FF70",X"FF82",X"FFC2",X"0039",X"00D4",X"018A",X"0271",X"0370",X"045D",X"051D",X"05B4",
		X"0636",X"06A9",X"06F5",X"0720",X"074D",X"0761",X"07A8",X"082F",X"08DC",X"0968",X"09E2",X"0A79",X"0AD6",X"0B2F",X"0B55",X"0B5A",
		X"0B26",X"0AD0",X"0A83",X"0A2C",X"09B6",X"095C",X"091E",X"090F",X"0919",X"0936",X"0950",X"0920",X"08EB",X"08B0",X"0870",X"0801",
		X"0758",X"06A1",X"05C4",X"04F5",X"042E",X"0358",X"0259",X"0147",X"0056",X"FF46",X"FE52",X"FD59",X"FC6C",X"FB7D",X"FA71",X"F96D",
		X"F866",X"F746",X"F609",X"F4EB",X"F3CE",X"F2B6",X"F1B4",X"F0ED",X"F032",X"EF85",X"EF00",X"EEB1",X"EE88",X"EE89",X"EEB3",X"EEDA",
		X"EF0F",X"EF23",X"EF2E",X"EF4C",X"EF74",X"EF9E",X"EFC3",X"EFCF",X"F008",X"F06A",X"F0D0",X"F167",X"F1F3",X"F283",X"F2F6",X"F380",
		X"F3F4",X"F47B",X"F4F1",X"F573",X"F60F",X"F693",X"F735",X"F7FB",X"F8C9",X"F9AB",X"FAB5",X"FBB6",X"FCD0",X"FDEA",X"FEF9",X"FFEE",
		X"00EF",X"01D2",X"0291",X"0358",X"0408",X"04A3",X"0541",X"05F8",X"068A",X"06F3",X"077A",X"07FE",X"0857",X"08CF",X"0935",X"0991",
		X"0A0A",X"0A66",X"0AEC",X"0B79",X"0BFF",X"0C63",X"0CD8",X"0D60",X"0E06",X"0EA2",X"0F2A",X"0F9B",X"1018",X"10AB",X"110B",X"1161",
		X"11BE",X"120F",X"122E",X"121B",X"1206",X"11EA",X"11A7",X"1173",X"112F",X"109D",X"100F",X"0F8A",X"0EF4",X"0E5D",X"0D99",X"0CB1",
		X"0BC8",X"0AD9",X"09FB",X"0908",X"0818",X"074A",X"0661",X"05B5",X"04E6",X"0419",X"033F",X"0247",X"0162",X"006E",X"FF84",X"FE87",
		X"FD99",X"FCD6",X"FC42",X"FBA9",X"FB1E",X"FAB4",X"FA4A",X"F9EC",X"F974",X"F901",X"F856",X"F7B2",X"F72A",X"F689",X"F5CE",X"F521",
		X"F492",X"F40E",X"F3B7",X"F36B",X"F325",X"F2CF",X"F283",X"F22F",X"F1D9",X"F182",X"F124",X"F0E9",X"F098",X"F04D",X"F01D",X"F003",
		X"F002",X"F00E",X"F047",X"F08A",X"F0CB",X"F112",X"F15E",X"F1C1",X"F21F",X"F276",X"F293",X"F28F",X"F297",X"F2A2",X"F2A3",X"F267",
		X"F21F",X"F1DF",X"F1D0",X"F1FC",X"F24A",X"F2AB",X"F342",X"F408",X"F524",X"F66E",X"F7B4",X"F8F7",X"FA17",X"FB48",X"FC9E",X"FDE1",
		X"FEFD",X"0001",X"010F",X"022E",X"0375",X"04EF",X"067F",X"0814",X"09C9",X"0B7C",X"0D17",X"0EB7",X"1010",X"111E",X"1216",X"12EB",
		X"137D",X"13B7",X"13EA",X"1441",X"149F",X"151A",X"15C6",X"1668",X"1700",X"179C",X"186C",X"191D",X"197E",X"19BC",X"19BA",X"198F",
		X"1940",X"18CD",X"1818",X"171D",X"161B",X"152B",X"1432",X"1341",X"1248",X"116B",X"108F",X"0F8E",X"0E98",X"0D73",X"0C2E",X"0AD3",
		X"0958",X"07E3",X"064E",X"04C0",X"0329",X"0193",X"003D",X"FEF6",X"FDD7",X"FCD3",X"FBDD",X"FB1A",X"FA6A",X"F9DA",X"F936",X"F8A6",
		X"F82F",X"F7BC",X"F73E",X"F6C0",X"F634",X"F585",X"F4DD",X"F425",X"F375",X"F2DF",X"F258",X"F1FA",X"F1A8",X"F160",X"F131",X"F105",
		X"F0EE",X"F0B8",X"F068",X"EFFC",X"EF83",X"EEED",X"EE5D",X"EE08",X"EDC3",X"ED79",X"ED31",X"ED21",X"ED2E",X"ED4D",X"ED84",X"EDC6",
		X"EE01",X"EE49",X"EE9D",X"EECE",X"EEF8",X"EEE3",X"EEB4",X"EE79",X"EE44",X"EE5F",X"EE62",X"EE88",X"EEB7",X"EF2B",X"EFCF",X"F070",
		X"F110",X"F17B",X"F1E0",X"F252",X"F2DF",X"F33D",X"F3B3",X"F429",X"F4FD",X"F5F6",X"F72E",X"F895",X"FA07",X"FB8F",X"FD17",X"FEBE",
		X"0029",X"0186",X"02F9",X"0435",X"0572",X"06B0",X"07C2",X"08F7",X"09FD",X"0B22",X"0C47",X"0D2E",X"0E13",X"0ECC",X"0F6A",X"0FFC",
		X"1054",X"10AB",X"10E9",X"1138",X"1172",X"1172",X"11A1",X"11E1",X"1257",X"12D3",X"1344",X"13C4",X"143B",X"1498",X"14D8",X"14F0",
		X"1509",X"14F7",X"14C4",X"148A",X"1461",X"1458",X"1434",X"1429",X"140D",X"13FC",X"13F2",X"1409",X"140D",X"13EA",X"138E",X"12F2",
		X"1248",X"118F",X"10BA",X"0FEF",X"0F09",X"0E23",X"0D4B",X"0C96",X"0BE2",X"0B64",X"0AF5",X"0A85",X"0A21",X"09A4",X"0914",X"0855",
		X"07A7",X"06E2",X"05F4",X"04E8",X"03DA",X"02BB",X"019D",X"008B",X"FF5B",X"FE2A",X"FCD6",X"FB7C",X"FA17",X"F89F",X"F73F",X"F5FA",
		X"F4AF",X"F355",X"F225",X"F117",X"F037",X"EF43",X"EE63",X"ED82",X"EC98",X"EBE1",X"EB3C",X"EACC",X"EA5E",X"E9FE",X"E9A6",X"E98F",
		X"E971",X"E959",X"E95B",X"E947",X"E92C",X"E8F6",X"E8DB",X"E8C0",X"E89D",X"E897",X"E8AA",X"E8BE",X"E90B",X"E966",X"E9EF",X"EA9B",
		X"EB66",X"EC42",X"ECFC",X"ED9E",X"EE6A",X"EF27",X"EFE2",X"F0A5",X"F147",X"F1E8",X"F2B1",X"F38F",X"F492",X"F577",X"F634",X"F71C",
		X"F7EB",X"F8D2",X"F9B6",X"FA65",X"FACE",X"FB31",X"FBB5",X"FC43",X"FCDC",X"FD65",X"FDDB",X"FE6B",X"FF32",X"003D",X"0160",X"0260",
		X"0351",X"0467",X"054E",X"0629",X"06F8",X"079C",X"0811",X"0869",X"08D1",X"092F",X"09AA",X"0A40",X"0AEE",X"0BAC",X"0C7B",X"0D8B",
		X"0E9C",X"0F9B",X"1086",X"113E",X"11F8",X"127A",X"12E7",X"133B",X"1369",X"13AB",X"1405",X"1462",X"14DB",X"1554",X"15E1",X"16A7",
		X"174A",X"17F7",X"186B",X"18CC",X"190C",X"1953",X"1972",X"1982",X"1966",X"1947",X"1929",X"18F3",X"189A",X"17EC",X"1751",X"16A8",
		X"15DF",X"14D5",X"13BF",X"129E",X"1191",X"106D",X"0F54",X"0E35",X"0D38",X"0C3D",X"0B33",X"0A20",X"0904",X"07B6",X"0646",X"04E2",
		X"0378",X"020B",X"0084",X"FF2F",X"FDCB",X"FC6E",X"FB2B",X"F9FC",X"F8B7",X"F775",X"F639",X"F4D4",X"F35D",X"F1F6",X"F085",X"EF2B",
		X"EDE8",X"ECBC",X"EBB7",X"EAC7",X"EA13",X"E980",X"E932",X"E8EF",X"E8B5",X"E865",X"E82C",X"E7E3",X"E789",X"E725",X"E69F",X"E62F",
		X"E5C3",X"E57C",X"E555",X"E565",X"E58F",X"E5C9",X"E61F",X"E69F",X"E726",X"E7B0",X"E814",X"E872",X"E8CF",X"E8EA",X"E90D",X"E91F",
		X"E94D",X"E998",X"E9F4",X"EA5D",X"EAF6",X"EBCF",X"ECFA",X"EE5D",X"EFD6",X"F165",X"F2F9",X"F48F",X"F60E",X"F781",X"F8C3",X"FA0B",
		X"FB24",X"FC4D",X"FD94",X"FEE8",X"004B",X"01B7",X"0344",X"04CC",X"0636",X"079D",X"0910",X"0A53",X"0B70",X"0C39",X"0CFF",X"0DAC",
		X"0E4A",X"0EEC",X"0FAB",X"106E",X"1127",X"120C",X"12F6",X"13CE",X"14A4",X"1541",X"15AD",X"15F8",X"161E",X"164E",X"1660",X"1679",
		X"1685",X"1699",X"16D0",X"1706",X"173D",X"177F",X"17C6",X"180C",X"182E",X"1803",X"17C7",X"176A",X"1706",X"167B",X"15CB",X"14E8",
		X"13F3",X"1309",X"1241",X"11B2",X"111E",X"108D",X"1006",X"0F93",X"0F4A",X"0F38",X"0F02",X"0ECD",X"0E6C",X"0DF3",X"0D57",X"0C9C",
		X"0BE2",X"0B17",X"0A42",X"0971",X"08B4",X"07F7",X"076E",X"06E5",X"0672",X"05FC",X"0590",X"0525",X"049E",X"0407",X"0348",X"028B",
		X"0193",X"005E",X"FF0A",X"FDC2",X"FC77",X"FB31",X"F9FF",X"F8C5",X"F789",X"F653",X"F520",X"F3FD",X"F2C8",X"F188",X"F02A",X"EECA",
		X"ED38",X"EBD9",X"EA9F",X"E944",X"E815",X"E6DD",X"E5CC",X"E4D1",X"E403",X"E38E",X"E348",X"E2E2",X"E2A9",X"E276",X"E281",X"E28C",
		X"E285",X"E287",X"E256",X"E25E",X"E28F",X"E2D3",X"E306",X"E35B",X"E3B9",X"E44B",X"E516",X"E611",X"E716",X"E7ED",X"E8FA",X"E9F7",
		X"EAD3",X"EBA5",X"EC6C",X"ED0D",X"EDA0",X"EE41",X"EF16",X"F011",X"F104",X"F231",X"F391",X"F51D",X"F6AB",X"F84B",X"FA11",X"FBBE",
		X"FD68",X"FF03",X"0078",X"01E4",X"031F",X"046D",X"05CD",X"073F",X"08C1",X"0A49",X"0BDE",X"0D77",X"0F21",X"10AB",X"11F6",X"131A",
		X"13E9",X"1498",X"152A",X"15AB",X"1624",X"1665",X"16C1",X"1726",X"17A9",X"1843",X"18CB",X"1961",X"1A04",X"1A9B",X"1B1B",X"1B93",
		X"1BE5",X"1C33",X"1C29",X"1C1F",X"1BF3",X"1B9E",X"1B28",X"1A8F",X"1A12",X"1986",X"1917",X"189A",X"1800",X"1776",X"16F1",X"166D",
		X"1609",X"1594",X"150A",X"1478",X"13E0",X"134B",X"128D",X"11D5",X"1119",X"1031",X"0F2B",X"0E17",X"0D17",X"0C15",X"0B02",X"09C6",
		X"0894",X"0765",X"0614",X"04E3",X"03CC",X"02A4",X"017E",X"0038",X"FF07",X"FDC0",X"FC83",X"FB64",X"FA33",X"F905",X"F7E6",X"F6CD",
		X"F5F0",X"F517",X"F45E",X"F3BA",X"F2EC",X"F24D",X"F19E",X"F101",X"F052",X"EFA6",X"EEE7",X"EE0D",X"ED55",X"ECB1",X"EBFE",X"EB44",
		X"EAB3",X"EA34",X"E9B9",X"E946",X"E8F2",X"E86D",X"E7F8",X"E78A",X"E6F4",X"E66A",X"E60B",X"E5C0",X"E57E",X"E53F",X"E502",X"E4EF",
		X"E52F",X"E5BE",X"E61A",X"E67E",X"E707",X"E768",X"E7E8",X"E861",X"E8CA",X"E92D",X"E987",X"EA05",X"EA95",X"EB56",X"EC30",X"ED22",
		X"EE06",X"EF17",X"F02B",X"F153",X"F265",X"F350",X"F438",X"F505",X"F5C0",X"F687",X"F763",X"F849",X"F971",X"FA9E",X"FBFB",X"FD7E",
		X"FF23",X"00C8",X"0292",X"0453",X"0620",X"07CC",X"0976",X"0B0E",X"0C71",X"0DE9",X"0F44",X"108A",X"1193",X"12AC",X"13C3",X"14CD",
		X"15D3",X"16C5",X"17AF",X"189C",X"197E",X"1A44",X"1B21",X"1BDC",X"1C6F",X"1CF0",X"1D73",X"1DE5",X"1E1F",X"1E1B",X"1E02",X"1DD3",
		X"1D92",X"1D27",X"1CA7",X"1C16",X"1B59",X"1AE1",X"1A90",X"1A2B",X"19BF",X"193F",X"18D9",X"1865",X"1800",X"17A4",X"170B",X"1658",
		X"157A",X"1491",X"13A6",X"12B8",X"11AA",X"1076",X"0F2B",X"0DDF",X"0C89",X"0B3D",X"0A05",X"08CB",X"0762",X"05F5",X"0490",X"034B",
		X"020B",X"00C5",X"FFB0",X"FE8E",X"FD76",X"FC57",X"FB4D",X"FA58",X"F98F",X"F8AC",X"F79F",X"F694",X"F584",X"F4C3",X"F3E7",X"F32F",
		X"F253",X"F18C",X"F0DA",X"F04E",X"EFD9",X"EF3B",X"EEA9",X"EE37",X"EDD0",X"ED5B",X"ECE9",X"EC6D",X"EBBE",X"EB13",X"EA79",X"E9CC",
		X"E941",X"E8A8",X"E816",X"E7A2",X"E75F",X"E734",X"E73C",X"E76D",X"E7C1",X"E80A",X"E859",X"E8C2",X"E925",X"E983",X"E9FB",X"EA90",
		X"EAF3",X"EB43",X"EBB4",X"EC24",X"ECA4",X"ED1B",X"ED86",X"EDE4",X"EE48",X"EEA9",X"EEE3",X"EF5F",X"EFD4",X"F05B",X"F102",X"F1A6",
		X"F249",X"F30C",X"F3ED",X"F4F6",X"F604",X"F715",X"F83D",X"F93A",X"FA38",X"FB36",X"FC50",X"FD6D",X"FE76",X"FF7E",X"00A9",X"01F0",
		X"034F",X"04A1",X"05D6",X"0708",X"0819",X"08FD",X"09CA",X"0A72",X"0AEB",X"0B26",X"0B56",X"0B90",X"0BCA",X"0C09",X"0C53",X"0CC2",
		X"0D45",X"0DF9",X"0E9B",X"0F3B",X"0FD7",X"1075",X"112B",X"11C4",X"124B",X"12B0",X"132B",X"1396",X"1418",X"14B1",X"1542",X"15BB",
		X"1639",X"16ED",X"177B",X"1800",X"1873",X"18C4",X"18E0",X"18F4",X"18FE",X"18CB",X"188F",X"1844",X"17F1",X"178A",X"1710",X"16CB",
		X"166F",X"15EA",X"154D",X"1497",X"13AD",X"1288",X"1177",X"1042",X"0F0B",X"0DCD",X"0C92",X"0B71",X"0A63",X"0966",X"087F",X"079B",
		X"06AB",X"05A0",X"0496",X"0392",X"0256",X"00FA",X"FF86",X"FE1A",X"FCAF",X"FB37",X"F9C9",X"F870",X"F72C",X"F60C",X"F512",X"F433",
		X"F34C",X"F276",X"F1AF",X"F103",X"F031",X"EF65",X"EEBE",X"EE01",X"ED5E",X"ECD4",X"EC60",X"EC09",X"EBCA",X"EBB7",X"EBB9",X"EBD3",
		X"EC15",X"EC45",X"EC75",X"ECAD",X"ECDA",X"ECEC",X"ED0A",X"ED19",X"ED14",X"ED09",X"ECF9",X"ED17",X"ED65",X"EDBE",X"EE47",X"EED8",
		X"EF6B",X"EFFF",X"F0C7",X"F17D",X"F208",X"F25F",X"F29A",X"F2C3",X"F2BC",X"F29A",X"F283",X"F299",X"F2B8",X"F2F4",X"F353",X"F3CC",
		X"F455",X"F4E5",X"F58D",X"F633",X"F6CB",X"F753",X"F7D8",X"F864",X"F8EF",X"F986",X"F9FB",X"FA78",X"FAFF",X"FBC2",X"FC9B",X"FD7C",
		X"FE58",X"FF3C",X"0016",X"00EB",X"01CB",X"02A1",X"0376",X"0436",X"04F4",X"05B8",X"065E",X"0700",X"078E",X"084E",X"090D",X"09E4",
		X"0AB0",X"0B7A",X"0C5B",X"0D12",X"0DB0",X"0E45",X"0EB3",X"0F10",X"0F69",X"0FB9",X"1010",X"1027",X"100E",X"0FD6",X"0FCB",X"0FA1",
		X"0F88",X"0F47",X"0F1B",X"0F0D",X"0F42",X"0F8A",X"0FD0",X"1023",X"106D",X"10B7",X"1106",X"1155",X"116A",X"1129",X"10BA",X"104A",
		X"0FF8",X"0FAA",X"0F4F",X"0EEE",X"0E99",X"0E6A",X"0E64",X"0E67",X"0E72",X"0E74",X"0E57",X"0E1D",X"0DE0",X"0D9D",X"0D3F",X"0CBB",
		X"0C0F",X"0B5C",X"0A99",X"09F0",X"0955",X"08D0",X"0834",X"0791",X"06CA",X"0613",X"0558",X"049A",X"03BA",X"02AF",X"0192",X"0088",
		X"FF5B",X"FE1D",X"FCDE",X"FB88",X"FA1C",X"F895",X"F72B",X"F5B0",X"F448",X"F2B2",X"F15B",X"F032",X"EF04",X"EE0E",X"ED45",X"EC92",
		X"EC00",X"EB9D",X"EB39",X"EAF3",X"EAAC",X"EA7F",X"EA4E",X"EA35",X"EA16",X"E9FF",X"E9EC",X"E9F4",X"EA10",X"EA0E",X"EA24",X"EA52",
		X"EA97",X"EABF",X"EAF4",X"EB3C",X"EB7C",X"EBBE",X"EC33",X"ECA8",X"ED43",X"EDFD",X"EEE0",X"F000",X"F11F",X"F24A",X"F38E",X"F4D3",
		X"F616",X"F776",X"F888",X"F97E",X"FA36",X"FACD",X"FB88",X"FC0C",X"FCCD",X"FD61",X"FE26",X"FEE4",X"FFAE",X"00A1",X"0193",X"02BE",
		X"03D4",X"04E8",X"05C0",X"0672",X"0717",X"078A",X"07F5",X"084B",X"0878",X"088C",X"08A4",X"08DF",X"0931",X"0997",X"0A1A",X"0AC8",
		X"0B61",X"0C39",X"0CE7",X"0DAB",X"0E4C",X"0E91",X"0EAE",X"0EA7",X"0EAD",X"0EA6",X"0EAB",X"0EAE",X"0E8D",X"0E53",X"0E48",X"0E54",
		X"0E75",X"0E92",X"0E8B",X"0E94",X"0E8E",X"0E98",X"0E9B",X"0EA5",X"0E8C",X"0E4D",X"0E26",X"0DE5",X"0DC6",X"0DA2",X"0D6C",X"0D29",
		X"0CB2",X"0C1F",X"0BA4",X"0B1B",X"0A82",X"09DB",X"0938",X"0894",X"07FF",X"078C",X"0718",X"06B1",X"065A",X"05BE",X"04EF",X"0435",
		X"036D",X"02A0",X"01CC",X"00ED",X"0022",X"FF5E",X"FEA2",X"FDF4",X"FD64",X"FCD2",X"FC50",X"FBD3",X"FB61",X"FAFA",X"FA5D",X"F9C9",
		X"F91A",X"F869",X"F7AF",X"F6FB",X"F67D",X"F608",X"F599",X"F549",X"F4E4",X"F492",X"F439",X"F3BE",X"F377",X"F34A",X"F31F",X"F2F1",
		X"F2CE",X"F291",X"F274",X"F258",X"F24F",X"F264",X"F277",X"F295",X"F2A3",X"F2D7",X"F313",X"F356",X"F397",X"F3D2",X"F40B",X"F418",
		X"F419",X"F429",X"F41B",X"F3FD",X"F3BF",X"F38A",X"F36B",X"F37E",X"F3B9",X"F405",X"F49B",X"F54E",X"F62E",X"F70B",X"F7EE",X"F8B6",
		X"F96E",X"F9E3",X"FA0E",X"FA0E",X"FA08",X"FA3E",X"FA6A",X"FAE6",X"FB85",X"FC4F",X"FD6E",X"FED7",X"0071",X"0228",X"03AF",X"04F4",
		X"0621",X"06FC",X"07CC",X"0882",X"0908",X"096F",X"09B6",X"0A09",X"0A99",X"0B76",X"0C6D",X"0D72",X"0E81",X"0F98",X"107E",X"117F",
		X"123F",X"12B6",X"12E4",X"12D1",X"12A9",X"123D",X"11CA",X"1148",X"10D5",X"1074",X"101D",X"0FEA",X"0FF2",X"0FDD",X"0FFD",X"1009",
		X"0FED",X"0FBD",X"0F74",X"0EE7",X"0E3D",X"0D82",X"0CB3",X"0BB7",X"0AA9",X"09A7",X"08AF",X"07D9",X"0727",X"066C",X"05B8",X"04EB",
		X"0436",X"037F",X"0289",X"0183",X"003E",X"FEEE",X"FD90",X"FC57",X"FB14",X"F9C3",X"F8A1",X"F7BE",X"F6FD",X"F675",X"F5FF",X"F5BA",
		X"F568",X"F520",X"F4EB",X"F4BB",X"F46C",X"F423",X"F3C3",X"F355",X"F2DC",X"F271",X"F210",X"F1AE",X"F1A7",X"F1CC",X"F220",X"F291",
		X"F301",X"F36B",X"F3D4",X"F44A",X"F4B5",X"F4DE",X"F4D8",X"F4C7",X"F48C",X"F44E",X"F425",X"F423",X"F441",X"F474",X"F508",X"F597",
		X"F63F",X"F708",X"F7D1",X"F89C",X"F92B",X"F9AC",X"FA27",X"FA7A",X"FAA1",X"FABC",X"FAEC",X"FAFE",X"FB15",X"FB43",X"FBA9",X"FC20",
		X"FCAE",X"FD3F",X"FDF4",X"FEA8",X"FF34",X"FFC3",X"0051",X"00D3",X"012C",X"018F",X"01E4",X"0236",X"029C",X"02F9",X"0370",X"03E3",
		X"0456",X"04C4",X"0511",X"055B",X"0594",X"05CE",X"0616",X"0679",X"06B7",X"06EA",X"071A",X"076F",X"079B",X"07D6",X"07FF",X"082E",
		X"085A",X"0851",X"0857",X"084D",X"0854",X"0830",X"07FA",X"07F2",X"07DB",X"07AC",X"079C",X"07B1",X"07B8",X"07C5",X"07D7",X"0808",
		X"0847",X"087F",X"08B0",X"08BF",X"08C7",X"08CA",X"08F0",X"08E0",X"08E8",X"08C8",X"0895",X"0852",X"07FB",X"07A1",X"0731",X"06B5",
		X"05FF",X"054E",X"04BB",X"0458",X"03F9",X"03AF",X"0371",X"0346",X"0344",X"0354",X"0377",X"0377",X"0367",X"0333",X"02E6",X"0293",
		X"020E",X"017E",X"00EF",X"0040",X"FFB5",X"FF46",X"FEE4",X"FEA2",X"FE50",X"FE0A",X"FDE5",X"FDC5",X"FD75",X"FD04",X"FC6C",X"FBA9",
		X"FAB1",X"F9B2",X"F8B4",X"F7BC",X"F6F5",X"F62F",X"F580",X"F4F1",X"F48F",X"F446",X"F423",X"F3FD",X"F402",X"F407",X"F411",X"F448",
		X"F461",X"F4A0",X"F4C2",X"F4E7",X"F522",X"F57B",X"F5EA",X"F644",X"F68C",X"F6D1",X"F723",X"F75F",X"F7AA",X"F807",X"F84A",X"F86C",
		X"F890",X"F8BE",X"F8F8",X"F94F",X"F9A6",X"FA08",X"FA65",X"FAF8",X"FBC4",X"FC93",X"FD7C",X"FE75",X"FF73",X"008D",X"01A5",X"02B6",
		X"03C9",X"04AD",X"0597",X"0688",X"0738",X"07B9",X"081F",X"0865",X"087B",X"0864",X"083A",X"07F9",X"07C4",X"078A",X"0753",X"0723",
		X"06E8",X"06D7",X"06EB",X"0701",X"0730",X"0778",X"07C1",X"081A",X"0880",X"08FB",X"0940",X"0977",X"0999",X"09C4",X"09E1",X"09DC",
		X"09D6",X"09C5",X"098F",X"0936",X"08C4",X"083E",X"07B0",X"070B",X"066F",X"0599",X"04B8",X"040B",X"0376",X"02D8",X"026F",X"0218",
		X"0191",X"0113",X"00AE",X"005E",X"0002",X"FF8F",X"FF3D",X"FED9",X"FEAB",X"FE8F",X"FE8D",X"FE77",X"FE53",X"FE3D",X"FE09",X"FDD2",
		X"FDB3",X"FD70",X"FD04",X"FC96",X"FC2A",X"FBB7",X"FB15",X"FA66",X"F9A2",X"F8D7",X"F823",X"F797",X"F711",X"F699",X"F62D",X"F5DC",
		X"F5C3",X"F592",X"F559",X"F540",X"F527",X"F534",X"F54A",X"F571",X"F5B9",X"F613",X"F689",X"F6FD",X"F789",X"F815",X"F890",X"F8FB",
		X"F963",X"F9E1",X"FA39",X"FA79",X"FABA",X"FB1E",X"FB7A",X"FBAF",X"FBDE",X"FC04",X"FC14",X"FC32",X"FC52",X"FC7B",X"FC8F",X"FC8E",
		X"FCA7",X"FCBC",X"FCD6",X"FD12",X"FD47",X"FD50",X"FD50",X"FD6C",X"FD8C",X"FDCB",X"FE00",X"FE3C",X"FE8B",X"FEB5",X"FF04",X"FF40",
		X"FF71",X"FF9D",X"FFC4",X"FFDB",X"FFE2",X"FFE8",X"FFF1",X"0009",X"0012",X"0001",X"FFE1",X"FFCE",X"FFDA",X"FFED",X"0045",X"00CE",
		X"0135",X"01D5",X"0287",X"033D",X"040E",X"04C3",X"056A",X"05E9",X"0670",X"0709",X"078A",X"080D",X"0898",X"0917",X"09C9",X"0A98",
		X"0B75",X"0C4A",X"0CFB",X"0DC9",X"0E8E",X"0F55",X"100F",X"1098",X"1105",X"1126",X"1125",X"1111",X"10E1",X"10A2",X"1075",X"1031",
		X"101D",X"0FEC",X"0FAA",X"0F70",X"0F29",X"0EDA",X"0E79",X"0DF8",X"0D48",X"0C7A",X"0B6D",X"0A5B",X"0905",X"07A7",X"0627",X"04A8",
		X"034B",X"020E",X"00FD",X"000D",X"FF3A",X"FE90",X"FE12",X"FDAD",X"FD39",X"FC9C",X"FBDF",X"FB2E",X"FA67",X"F9C1",X"F908",X"F83B",
		X"F78C",X"F6FA",X"F68C",X"F65A",X"F62B",X"F5FD",X"F5DE",X"F5B4",X"F595",X"F581",X"F554",X"F4FB",X"F496",X"F442",X"F3E9",X"F39B",
		X"F360",X"F341",X"F368",X"F3B5",X"F42B",X"F4AB",X"F51A",X"F581",X"F5DB",X"F634",X"F670",X"F691",X"F6BE",X"F6ED",X"F73C",X"F799",
		X"F80F",X"F852",X"F8CC",X"F92D",X"F97B",X"F9A8",X"F9AC",X"F96F",X"F928",X"F8EA",X"F8B9",X"F87F",X"F82E",X"F830",X"F83D",X"F876",
		X"F8C7",X"F900",X"F941",X"F981",X"F9EB",X"FA6A",X"FAD4",X"FB3C",X"FBB1",X"FC39",X"FD03",X"FDB8",X"FE65",X"FF0B",X"FF9F",X"0083",
		X"0138",X"020F",X"02C6",X"035C",X"03F8",X"047C",X"0505",X"0584",X"05E9",X"062D",X"0671",X"06A1",X"06C4",X"06D7",X"0718",X"0772",
		X"07BA",X"080B",X"0856",X"08B6",X"0929",X"09DA",X"0A82",X"0B28",X"0BB3",X"0C27",X"0CA0",X"0D05",X"0D7A",X"0DC7",X"0DDD",X"0DE2",
		X"0DDA",X"0DAD",X"0D74",X"0D0A",X"0C7F",X"0BBF",X"0AD1",X"09EE",X"08E7",X"07FF",X"0719",X"066C",X"05B2",X"0519",X"0498",X"0427",
		X"03CB",X"036B",X"0339",X"02EF",X"02C1",X"0275",X"022E",X"01DA",X"01B3",X"0188",X"0182",X"0188",X"01A5",X"01E0",X"01FF",X"0216",
		X"020C",X"01FF",X"01C0",X"0169",X"00DC",X"0038",X"FF9E",X"FF06",X"FE76",X"FDE0",X"FD52",X"FCD4",X"FC48",X"FBC1",X"FB27",X"FA7E",
		X"F9DF",X"F939",X"F88F",X"F806",X"F77E",X"F705",X"F6A5",X"F628",X"F5BA",X"F561",X"F514",X"F4DD",X"F4A8",X"F45A",X"F3F5",X"F39F",
		X"F348",X"F2EA",X"F28E",X"F217",X"F1C1",X"F175",X"F156",X"F138",X"F130",X"F140",X"F15A",X"F15A",X"F16C",X"F168",X"F139",X"F10A",
		X"F0BD",X"F081",X"F04A",X"F02F",X"F05E",X"F0B7",X"F136",X"F1E3",X"F2BA",X"F3C4",X"F50A",X"F66C",X"F79E",X"F8C3",X"F9F5",X"FB21",
		X"FC4B",X"FD74",X"FE64",X"FF50",X"0021",X"011D",X"0217",X"031E",X"0435",X"0535",X"0624",X"0716",X"0802",X"08F3",X"09DE",X"0AA1",
		X"0B4B",X"0BDD",X"0C46",X"0CC3",X"0D44",X"0DAF",X"0E14",X"0E7B",X"0ED7",X"0F3B",X"0FB0",X"1028",X"108A",X"10DF",X"1126",X"115B",
		X"11B1",X"11F4",X"1244",X"1283",X"12B2",X"12AD",X"1298",X"1289",X"127A",X"125D",X"1228",X"11C7",X"1157",X"10CF",X"102E",X"0F83",
		X"0EDC",X"0E2C",X"0D5E",X"0C82",X"0BB1",X"0ADA",X"09E0",X"08F6",X"0816",X"073B",X"064E",X"056C",X"04BD",X"0415",X"037F",X"02DD",
		X"025E",X"01CD",X"0144",X"00D6",X"0048",X"FFC9",X"FF3B",X"FEA6",X"FE0A",X"FD38",X"FC80",X"FBE2",X"FB41",X"FAAB",X"FA14",X"F957",
		X"F89D",X"F809",X"F766",X"F6B9",X"F634",X"F5CD",X"F53F",X"F4B8",X"F454",X"F418",X"F3F8",X"F3ED",X"F3C3",X"F38C",X"F367",X"F31D",
		X"F2DD",X"F29C",X"F23F",X"F1D7",X"F168",X"F12D",X"F10E",X"F134",X"F16E",X"F1A1",X"F1EB",X"F23E",X"F2D2",X"F38F",X"F444",X"F4F4",
		X"F55B",X"F5A0",X"F5DD",X"F619",X"F66B",X"F69B",X"F6D1",X"F70B",X"F761",X"F7F7",X"F87A",X"F928",X"F9BC",X"FA39",X"FAC2",X"FB39",
		X"FBCB",X"FC56",X"FCDE",X"FD55",X"FDE9",X"FE7D",X"FF0F",X"FFBC",X"006F",X"010C",X"01A9",X"0242",X"02CC",X"0347",X"038D",X"03AB",
		X"03B5",X"03A9",X"0398",X"0390",X"0381",X"0392",X"03E5",X"0448",X"04B4",X"052A",X"05BF",X"066A",X"070E",X"07A7",X"080D",X"0851",
		X"0896",X"08E2",X"091F",X"0950",X"0968",X"096A",X"0977",X"09A6",X"09EC",X"0A29",X"0A66",X"0AAA",X"0B01",X"0B57",X"0B90",X"0BDC",
		X"0C0A",X"0C14",X"0BF7",X"0B98",X"0B10",X"0A3B",X"0972",X"0874",X"0792",X"06B2",X"05E4",X"055B",X"0518",X"0506",X"0506",X"0521",
		X"0553",X"0576",X"058D",X"0597",X"054B",X"04C6",X"03F9",X"02F3",X"01F1",X"0118",X"0048",X"FFAB",X"FF10",X"FEC1",X"FEAE",X"FEBD",
		X"FEC4",X"FED3",X"FEB3",X"FE6F",X"FE35",X"FDCA",X"FD45",X"FCBD",X"FC39",X"FBA6",X"FB42",X"FB05",X"FAE1",X"FAE9",X"FB27",X"FB76",
		X"FBC0",X"FBE8",X"FC0B",X"FC2C",X"FC3E",X"FC55",X"FC4D",X"FC20",X"FBE2",X"FBAE",X"FB82",X"FB46",X"FAF3",X"FAA1",X"FA8F",X"FA79",
		X"FA71",X"FA46",X"FA11",X"FA08",X"F9EC",X"F9DE",X"F9B9",X"F98E",X"F95E",X"F939",X"F90A",X"F8DC",X"F89C",X"F87E",X"F893",X"F8CE",
		X"F8E5",X"F8EB",X"F8ED",X"F8EF",X"F919",X"F942",X"F979",X"F983",X"F9BC",X"F9D7",X"F9E0",X"FA03",X"FA16",X"FA28",X"FA34",X"FA69",
		X"FAB0",X"FB1F",X"FBC0",X"FC56",X"FCE7",X"FD87",X"FE2C",X"FEDA",X"FF8D",X"0011",X"0074",X"00B2",X"00F2",X"0120",X"0142",X"0160",
		X"0171",X"01AB",X"01F4",X"024C",X"02B2",X"0310",X"0384",X"03FF",X"0470",X"04D3",X"04FF",X"050F",X"0528",X"0541",X"0535",X"0504",
		X"04CB",X"0496",X"0462",X"0452",X"045D",X"0467",X"0466",X"0465",X"0469",X"0463",X"047B",X"048F",X"048E",X"048A",X"0485",X"0485",
		X"048A",X"0482",X"0478",X"046A",X"0442",X"040C",X"03B4",X"0358",X"02F8",X"02AB",X"02A0",X"025C",X"0227",X"0215",X"0201",X"01FB",
		X"01F0",X"01CA",X"019D",X"016C",X"0168",X"0157",X"0168",X"0192",X"01AD",X"01CF",X"021C",X"028E",X"031B",X"03B3",X"044F",X"04D7",
		X"0541",X"05B0",X"0615",X"0669",X"066C",X"065D",X"0626",X"05EF",X"05AE",X"057C",X"054E",X"0510",X"04D1",X"04B9",X"049A",X"044F",
		X"03F8",X"0393",X"0336",X"02A4",X"01EC",X"0142",X"0080",X"FFE1",X"FF53",X"FEB2",X"FE2E",X"FDA0",X"FD4A",X"FD46",X"FD1C",X"FCDB",
		X"FC9A",X"FC4E",X"FBF6",X"FB8A",X"FB1C",X"FAA2",X"F9E6",X"F95C",X"F8D7",X"F857",X"F805",X"F7A4",X"F76B",X"F737",X"F708",X"F6CC",
		X"F698",X"F67A",X"F65D",X"F621",X"F5FA",X"F5D9",X"F5EA",X"F613",X"F619",X"F622",X"F620",X"F614",X"F606",X"F5FB",X"F601",X"F603",
		X"F61F",X"F667",X"F6C7",X"F773",X"F855",X"F95C",X"FA68",X"FB5B",X"FC5B",X"FD39",X"FE23",X"FEDC",X"FF28",X"FF43",X"FF06",X"FEEE",
		X"FEDD",X"FF04",X"FF48",X"FFB9",X"0060",X"012B",X"0207",X"02EA",X"03F4",X"04D0",X"0598",X"05FE",X"0656",X"0696",X"06BA",X"06ED",
		X"0723",X"076D",X"07C7",X"0838",X"08DD",X"09A9",X"0A53",X"0ABD",X"0AEC",X"0B21",X"0B48",X"0B09",X"0AB0",X"0A42",X"09A9",X"094F",
		X"091D",X"090E",X"08FE",X"0907",X"091A",X"0920",X"0937",X"0953",X"0948",X"090B",X"08B0",X"083E",X"07AE",X"0712",X"06A0",X"062D",
		X"0598",X"04F6",X"0493",X"041A",X"03CF",X"03A9",X"0384",X"0340",X"0305",X"02BA",X"0273",X"0247",X"021E",X"01EA",X"0192",X"0144",
		X"00F1",X"00C2",X"0092",X"005E",X"001B",X"FFC0",X"FF86",X"FF48",X"FEFF",X"FEB8",X"FE51",X"FE00",X"FDB1",X"FD77",X"FD33",X"FD0F",
		X"FCC5",X"FC8A",X"FC32",X"FBD2",X"FB62",X"FADA",X"FA50",X"F9B3",X"F8ED",X"F851",X"F7CA",X"F728",X"F6DC",X"F673",X"F639",X"F628",
		X"F625",X"F605",X"F5EC",X"F5DF",X"F5B0",X"F578",X"F522",X"F4CF",X"F475",X"F41E",X"F3F5",X"F3CB",X"F383",X"F359",X"F33A",X"F349",
		X"F388",X"F3CC",X"F3E2",X"F3DF",X"F3C9",X"F3CF",X"F40C",X"F44C",X"F482",X"F4A1",X"F4E2",X"F53F",X"F5EA",X"F687",X"F749",X"F7EC",
		X"F888",X"F93C",X"FA02",X"FAFF",X"FBDC",X"FCBD",X"FD98",X"FE74",X"FF42",X"0016",X"00DE",X"01C8",X"02A0",X"034A",X"03D7",X"0468",
		X"0525",X"05D4",X"06B2",X"0761",X"07F9",X"0891",X"093A",X"09DB",X"0A82",X"0B2A",X"0B76",X"0BC7",X"0C00",X"0C6E",X"0CBA",X"0CF3",
		X"0D0E",X"0D0C",X"0D19",X"0D49",X"0D96",X"0DC6",X"0DF9",X"0E09",X"0DEE",X"0DC7",X"0DA9",X"0D79",X"0D4A",X"0CEB",X"0C83",X"0C23",
		X"0B8E",X"0B1A",X"0AF1",X"0AD7",X"0A9C",X"0A4C",X"0A0B",X"09AE",X"095E",X"0910",X"0881",X"07D1",X"06FF",X"0640",X"05B6",X"0558",
		X"0520",X"04CD",X"0490",X"0475",X"0467",X"044E",X"0435",X"03DE",X"036D",X"02F7",X"0285",X"020B",X"016A",X"00C9",X"0022",X"FF88",
		X"FF23",X"FEE9",X"FE90",X"FE25",X"FDAE",X"FD5F",X"FCED",X"FC81",X"FC11",X"FB96",X"FB00",X"FA70",X"F9EC",X"F989",X"F913",X"F8B6",
		X"F87C",X"F832",X"F7E6",X"F799",X"F784",X"F781",X"F77A",X"F722",X"F6E4",X"F6AC",X"F68A",X"F68C",X"F666",X"F633",X"F60D",X"F611",
		X"F638",X"F665",X"F690",X"F6B7",X"F6CB",X"F6EC",X"F6FC",X"F70C",X"F72C",X"F744",X"F733",X"F716",X"F723",X"F750",X"F770",X"F7BE",
		X"F811",X"F847",X"F893",X"F8FC",X"F96C",X"F9C8",X"F9F6",X"FA03",X"FA28",X"FA75",X"FADC",X"FB3E",X"FB97",X"FBF5",X"FC5A",X"FCC7",
		X"FD40",X"FDD0",X"FE59",X"FEB7",X"FEF3",X"FF24",X"FF64",X"FF8C",X"FFA9",X"FFB2",X"FFAC",X"FFAE",X"FFDF",X"002A",X"0088",X"00F0",
		X"0143",X"0199",X"01F6",X"0264",X"02D5",X"0347",X"0398",X"03CA",X"03F0",X"0419",X"043F",X"045F",X"048D",X"0489",X"04B6",X"04BB",
		X"049F",X"0483",X"0454",X"040A",X"0398",X"0330",X"02F5",X"02E1",X"02F8",X"0340",X"03AC",X"044D",X"04FC",X"05C5",X"06B5",X"077A",
		X"080D",X"0863",X"08B0",X"08C4",X"08B0",X"08BB",X"0897",X"08B2",X"08B6",X"08C2",X"08DD",X"08FE",X"0931",X"095F",X"0977",X"09B5",
		X"09E7",X"09F7",X"0A10",X"09CF",X"0967",X"08EA",X"0861",X"07BF",X"072F",X"0689",X"05CA",X"04EE",X"0434",X"03B9",X"036E",X"0349",
		X"032A",X"0341",X"0380",X"03CD",X"0426",X"0448",X"0436",X"0405",X"03CC",X"0351",X"028C",X"0199",X"0078",X"FF6A",X"FE75",X"FDB6",
		X"FCE3",X"FC3A",X"FBA9",X"FAFC",X"FA80",X"F9F8",X"F98E",X"F92A",X"F8E2",X"F8A3",X"F85C",X"F835",X"F7DA",X"F7A7",X"F772",X"F771",
		X"F790",X"F7DF",X"F82E",X"F87D",X"F8CB",X"F904",X"F941",X"F967",X"F991",X"F9C4",X"F9F2",X"FA01",X"F9F1",X"F9F9",X"F9E8",X"FA07",
		X"FA3A",X"FA54",X"FA51",X"FA7C",X"FA99",X"FAAD",X"FAB9",X"FA75",X"F9F8",X"F942",X"F8A3",X"F815",X"F788",X"F71F",X"F6A2",X"F646",
		X"F61C",X"F610",X"F661",X"F6B7",X"F732",X"F7A9",X"F817",X"F85D",X"F898",X"F8E7",X"F913",X"F91A",X"F90C",X"F8F5",X"F8CB",X"F8C7",
		X"F8FC",X"F934",X"F973",X"F9C0",X"FA20",X"FA8E",X"FB2A",X"FBA9",X"FC3A",X"FCB6",X"FD3E",X"FDA8",X"FE21",X"FE8A",X"FEFC",X"FF64",
		X"FFC8",X"0058",X"00E2",X"0183",X"0219",X"02C1",X"034B",X"03F6",X"04A7",X"054E",X"05E0",X"0636",X"0677",X"0686",X"069C",X"06CF",
		X"0705",X"0763",X"07C0",X"0832",X"08B5",X"0960",X"0A43",X"0B2D",X"0BFE",X"0CC1",X"0D4B",X"0DE9",X"0E60",X"0ED4",X"0F2C",X"0F51",
		X"0F53",X"0F5E",X"0F64",X"0F52",X"0F48",X"0F2E",X"0F13",X"0ED8",X"0EA7",X"0EA1",X"0E9D",X"0EC6",X"0ED5",X"0EF4",X"0F11",X"0F29",
		X"0F4B",X"0F4F",X"0F33",X"0EFF",X"0EB5",X"0E3C",X"0DD5",X"0D52",X"0CCD",X"0C1A",X"0B62",X"0AB6",X"09F9",X"0933",X"0882",X"07D5",
		X"06F3",X"0605",X"0519",X"0419",X"0317",X"01FD",X"00E6",X"FFBB",X"FEA1",X"FD92",X"FC78",X"FB7C",X"FA82",X"F9A2",X"F8A5",X"F7B3",
		X"F6CF",X"F5E8",X"F518",X"F451",X"F393",X"F2CF",X"F241",X"F1A7",X"F119",X"F0CB",X"F089",X"F062",X"F050",X"F048",X"F040",X"F02D",
		X"F038",X"F032",X"F01D",X"EFF2",X"EFB3",X"EF83",X"EF49",X"EF03",X"EED2",X"EE9B",X"EE69",X"EE50",X"EE7D",X"EEE1",X"EF62",X"EFF3",
		X"F075",X"F0EC",X"F187",X"F215",X"F2B5",X"F318",X"F37C",X"F3A6",X"F3CB",X"F403",X"F410",X"F430",X"F42D",X"F430",X"F426",X"F41C",
		X"F40A",X"F3FF",X"F409",X"F432",X"F430",X"F440",X"F460",X"F4B6",X"F529",X"F5AF",X"F67F",X"F763",X"F867",X"F995",X"FAAF",X"FBE8",
		X"FD2E",X"FE3D",X"FF64",X"0057",X"015D",X"0240",X"031F",X"0402",X"04AD",X"0580",X"065D",X"075B",X"085A",X"096D",X"0A7C",X"0B9E",
		X"0CD7",X"0E04",X"0F2F",X"105B",X"118C",X"12C4",X"13EB",X"1502",X"160C",X"16CC",X"1767",X"17F9",X"1887",X"18ED",X"192A",X"1967",
		X"198D",X"199C",X"198E",X"198D",X"1969",X"1943",X"18FE",X"18CE",X"187B",X"1816",X"17BB",X"170F",X"1646",X"155A",X"145A",X"1326",
		X"11C5",X"1057",X"0EC3",X"0D46",X"0BEA",X"0AA9",X"09A8",X"08E9",X"085C",X"07DE",X"075F",X"06DE",X"0673",X"05E2",X"053D",X"0454",
		X"0344",X"0210",X"00D3",X"FF92",X"FE5B",X"FD3D",X"FC38",X"FB29",X"FA45",X"F99D",X"F900",X"F87D",X"F7E5",X"F72F",X"F64B",X"F574",
		X"F479",X"F377",X"F274",X"F177",X"F08A",X"EFC8",X"EF67",X"EF22",X"EEFC",X"EEDE",X"EEBE",X"EE94",X"EE45",X"EDFD",X"ED84",X"ECF6",
		X"EC57",X"EBCD",X"EB40",X"EA97",X"EA15",X"E9C0",X"E975",X"E94E",X"E92C",X"E93D",X"E957",X"E9AC",X"E9EA",X"EA25",X"EA5B",X"EAB6",
		X"EB23",X"EB9E",X"EC26",X"ECB2",X"ED4C",X"EDB6",X"EE5F",X"EEF9",X"EFC3",X"F076",X"F12B",X"F1CD",X"F28D",X"F339",X"F3F5",X"F4B7",
		X"F5B3",X"F6B7",X"F7E8",X"F951",X"FAB7",X"FC42",X"FDDA",X"FF5C",X"00A9",X"01E8",X"0326",X"0449",X"0534",X"0625",X"06EE",X"07C8",
		X"08F2",X"0A2A",X"0B68",X"0CBE",X"0E29",X"0F6F",X"10D1",X"122C",X"133E",X"1409",X"1499",X"1510",X"1582",X"15F4",X"1646",X"1664",
		X"167E",X"1696",X"16F4",X"175F",X"17B3",X"17FB",X"1813",X"17F1",X"179E",X"1736",X"16A4",X"15C1",X"14D1",X"13EF",X"12EB",X"1234",
		X"11C9",X"116A",X"112F",X"10EF",X"10BB",X"10A1",X"1074",X"1049",X"0FDD",X"0F2C",X"0E41",X"0D30",X"0C24",X"0B0D",X"09EF",X"08C6",
		X"0792",X"0682",X"05B9",X"0534",X"04DD",X"0494",X"043E",X"03D8",X"037D",X"0359",X"0318",X"02C0",X"01FF",X"00FF",X"FFDF",X"FEC7",
		X"FDAC",X"FCBA",X"FBB6",X"FAB3",X"F9B0",X"F8E1",X"F85D",X"F80E",X"F7F1",X"F7D1",X"F771",X"F6EC",X"F63A",X"F552",X"F451",X"F32B",
		X"F1D6",X"F041",X"EEBD",X"ED61",X"EC5C",X"EBA4",X"EB4E",X"EB3D",X"EB31",X"EB61",X"EBD4",X"EC3D",X"EC7D",X"EC78",X"EC4C",X"EBDD",
		X"EB57",X"EABA",X"EA34",X"E9C4",X"E99A",X"E99D",X"E9DF",X"EA71",X"EB2E",X"EC48",X"ED5C",X"EE61",X"EF4B",X"F02C",X"F0D5",X"F151",
		X"F193",X"F1B9",X"F1E0",X"F230",X"F2C7",X"F380",X"F483",X"F5AE",X"F705",X"F867",X"F9C2",X"FB18",X"FC4D",X"FD61",X"FE3D",X"FED2",
		X"FF62",X"FFD0",X"0068",X"010B",X"01A3",X"0258",X"034D",X"0423",X"04FB",X"05E9",X"06C9",X"078B",X"081E",X"0893",X"090C",X"096A",
		X"09B4",X"09E8",X"09EA",X"09F4",X"0A1F",X"0A7C",X"0AF7",X"0B6C",X"0BDE",X"0C71",X"0CE6",X"0D75",X"0DEE",X"0E57",X"0EB2",X"0F11",
		X"0F55",X"0F82",X"0F93",X"0F99",X"0F8D",X"0F3C",X"0EDB",X"0E6B",X"0DEC",X"0D4B",X"0CE3",X"0CAE",X"0C7D",X"0C82",X"0CA2",X"0CDB",
		X"0D64",X"0E06",X"0EA2",X"0F0E",X"0F38",X"0F42",X"0F53",X"0F52",X"0F35",X"0F25",X"0F12",X"0EE1",X"0EC0",X"0EEB",X"0EF5",X"0F06",
		X"0F12",X"0F01",X"0EB4",X"0E5F",X"0DD9",X"0D28",X"0C77",X"0B9A",X"0AA8",X"09B9",X"08A7",X"07B7",X"06D1",X"05EC",X"0550",X"048C",
		X"03E2",X"031D",X"0244",X"016E",X"005A",X"FF37",X"FE28",X"FD1A",X"FC33",X"FB41",X"FA56",X"F98A",X"F8C8",X"F839",X"F79F",X"F719",
		X"F694",X"F5F5",X"F530",X"F452",X"F39E",X"F2DC",X"F20B",X"F14C",X"F071",X"EF90",X"EEDD",X"EE52",X"EDF7",X"ED8B",X"ECF8",X"EC6A",
		X"EBC8",X"EB32",X"EAB3",X"EA50",X"E9B6",X"E918",X"E876",X"E7EF",X"E79F",X"E79E",X"E7CA",X"E7E7",X"E80A",X"E849",X"E8D2",X"E96E",
		X"EA1F",X"EADB",X"EB91",X"EC39",X"ECDF",X"EDB8",X"EE88",X"EF74",X"F073",X"F181",X"F27A",X"F37E",X"F497",X"F5B0",X"F6F9",X"F80A",
		X"F8F6",X"F9FC",X"FAFE",X"FC04",X"FCE6",X"FDAA",X"FE71",X"FEEA",X"FF63",X"FFD1",X"0054",X"00C8",X"0153",X"01F0",X"029A",X"0370",
		X"044C",X"0537",X"0618",X"072E",X"084C",X"094A",X"0A32",X"0B02",X"0BBC",X"0C64",X"0D23",X"0DCD",X"0E68",X"0EF9",X"0F76",X"100D",
		X"10B0",X"113F",X"11BA",X"11F2",X"11F7",X"11DB",X"119A",X"1158",X"10F3",X"1065",X"0FD4",X"0F33",X"0ED1",X"0E93",X"0E8C",X"0EC3",
		X"0EF4",X"0F4F",X"0FB5",X"102D",X"1092",X"10EE",X"1117",X"1113",X"10E9",X"10C8",X"1081",X"1042",X"100E",X"0FDF",X"0FE1",X"0FE2",
		X"1008",X"1028",X"1033",X"1013",X"0FDF",X"0F71",X"0EE5",X"0E1F",X"0D23",X"0C12",X"0ADC",X"09AC",X"0863",X"0712",X"05F5",X"04EB",
		X"040D",X"0322",X"0269",X"01BF",X"0137",X"00BC",X"0022",X"FF77",X"FEA5",X"FDC0",X"FCE1",X"FC10",X"FB3B",X"FA53",X"F947",X"F842",
		X"F763",X"F691",X"F5C3",X"F536",X"F497",X"F3EE",X"F344",X"F292",X"F211",X"F18C",X"F0EC",X"F033",X"EF49",X"EE80",X"EDE4",X"ED53",
		X"ECA5",X"EC0B",X"EB79",X"EB03",X"EAAD",X"EA80",X"EA6B",X"EA69",X"EA56",X"EA56",X"EA57",X"EA7C",X"EAB1",X"EAFA",X"EB74",X"EC07",
		X"ECB3",X"ED72",X"EE66",X"EF62",X"F07F",X"F16A",X"F26C",X"F33A",X"F410",X"F4DE",X"F579",X"F620",X"F698",X"F709",X"F765",X"F7CB",
		X"F871",X"F93A",X"FA07",X"FACD",X"FB79",X"FC0B",X"FCB1",X"FD61",X"FE1B",X"FE99",X"FEF9",X"FF5D",X"FF9C",X"FFDE",X"0037",X"00AF",
		X"011A",X"01CB",X"0290",X"0356",X"045F",X"0581",X"06D2",X"0819",X"0949",X"0A6B",X"0B3D",X"0BF1",X"0C87",X"0CED",X"0D2C",X"0D2A",
		X"0D27",X"0D32",X"0D3B",X"0D6F",X"0DE1",X"0E4B",X"0EB7",X"0F17",X"0F69",X"0FC1",X"1012",X"104E",X"1045",X"1010",X"0FCF",X"0F95",
		X"0F58",X"0F28",X"0EE5",X"0EAA",X"0E84",X"0E89",X"0E88",X"0E9B",X"0EBC",X"0EB6",X"0EA7",X"0E87",X"0E6A",X"0E18",X"0D8F",X"0CFB",
		X"0C6E",X"0BA8",X"0AF4",X"0A5A",X"09E3",X"095D",X"08B6",X"0832",X"07D0",X"0782",X"0724",X"068B",X"05A1",X"0499",X"0387",X"025E",
		X"013D",X"FFE5",X"FE83",X"FD42",X"FC2D",X"FB4D",X"FAAE",X"FA37",X"F9EF",X"F9CE",X"F9CE",X"F9CD",X"F9DB",X"F9C7",X"F985",X"F935",
		X"F8D9",X"F85C",X"F7B7",X"F71B",X"F6AE",X"F648",X"F602",X"F5FD",X"F5F7",X"F613",X"F624",X"F669",X"F6DA",X"F718",X"F74D",X"F772",
		X"F777",X"F798",X"F7BF",X"F7F3",X"F802",X"F81B",X"F83C",X"F864",X"F88E",X"F8CD",X"F905",X"F928",X"F932",X"F951",X"F999",X"F9E4",
		X"FA10",X"FA37",X"FA3F",X"FA29",X"F9FD",X"F9AB",X"F95E",X"F8E9",X"F887",X"F843",X"F801",X"F7E4",X"F7F7",X"F82F",X"F88A",X"F8C9",
		X"F8E7",X"F8F1",X"F8C8",X"F87D",X"F82D",X"F7D5",X"F77C",X"F6FB",X"F6A3",X"F66E",X"F67B",X"F702",X"F7CC",X"F8C3",X"F9A9",X"FAB5",
		X"FBDD",X"FCFC",X"FE02",X"FED2",X"FF59",X"FF94",X"FFCF",X"0020",X"0075",X"00AB",X"00F7",X"0140",X"0191",X"0213",X"028D",X"0320",
		X"03B5",X"043A",X"04CE",X"0543",X"05CA",X"0657",X"06DC",X"0774",X"07F9",X"085E",X"08A0",X"090D",X"0985",X"09F9",X"0A4C",X"0A89",
		X"0AA3",X"0AAB",X"0AE6",X"0B22",X"0B2B",X"0AF6",X"0ACA",X"0A76",X"0A15",X"09F5",X"09D9",X"098B",X"0958",X"092B",X"0904",X"0907",
		X"0925",X"0930",X"0941",X"093D",X"093F",X"0955",X"0966",X"0965",X"092F",X"08BF",X"0856",X"07FA",X"077A",X"06D8",X"063D",X"05B4",
		X"052A",X"049E",X"041A",X"03AB",X"0344",X"0328",X"0305",X"02FB",X"02D5",X"02A6",X"026E",X"0231",X"01EE",X"0162",X"00D0",X"0019",
		X"FF82",X"FF19",X"FEB9",X"FE4A",X"FDFD",X"FDC9",X"FDA7",X"FD87",X"FD60",X"FD3C",X"FD05",X"FC96",X"FBF5",X"FB61",X"FABE",X"FA25",
		X"F998",X"F916",X"F8BA",X"F862",X"F858",X"F873",X"F898",X"F89D",X"F876",X"F836",X"F7E0",X"F785",X"F730",X"F6F5",X"F6C2",X"F6D1",
		X"F6F5",X"F731",X"F79C",X"F811",X"F887",X"F90D",X"F990",X"F9DC",X"FA01",X"FA24",X"FA03",X"F9B9",X"F966",X"F8F1",X"F860",X"F80B",
		X"F7DB",X"F7C1",X"F78E",X"F783",X"F77B",X"F76F",X"F79E",X"F7DC",X"F80F",X"F827",X"F845",X"F83F",X"F83F",X"F83E",X"F843",X"F848",
		X"F83B",X"F841",X"F849",X"F89D",X"F907",X"F995",X"FA2E",X"FAB3",X"FB74",X"FC73",X"FDA3",X"FEBD",X"FFE3",X"0110",X"020E",X"031C",
		X"042A",X"0543",X"064A",X"071F",X"07E5",X"087E",X"090F",X"098B",X"09EB",X"0A39",X"0A7B",X"0AB9",X"0AF4",X"0B50",X"0BB2",X"0C3C",
		X"0CD8",X"0D4F",X"0DD1",X"0E3C",X"0E9C",X"0EC8",X"0EDC",X"0ECE",X"0EB3",X"0EAA",X"0E88",X"0E68",X"0E2C",X"0DF1",X"0DA5",X"0D96",
		X"0D8F",X"0D66",X"0D48",X"0D01",X"0CA5",X"0C22",X"0BD4",X"0B51",X"0AC1",X"0A04",X"0928",X"0856",X"07A1",X"06FC",X"0617",X"0556",
		X"0489",X"03AE",X"02D6",X"022C",X"01AA",X"0113",X"0078",X"FFF9",X"FF8D",X"FF0E",X"FE82",X"FE1C",X"FD95",X"FCF5",X"FC51",X"FB8E",
		X"FAE4",X"FA38",X"F99C",X"F932",X"F8BF",X"F853",X"F7FE",X"F7C2",X"F794",X"F750",X"F6F0",X"F668",X"F5C7",X"F511",X"F435",X"F35C",
		X"F276",X"F1C2",X"F119",X"F077",X"F01B",X"EFFD",X"F01B",X"F03A",X"F050",X"F060",X"F066",X"F06F",X"F07A",X"F08D",X"F0A1",X"F0BD",
		X"F0C5",X"F102",X"F17D",X"F21D",X"F2FC",X"F3D1",X"F4BF",X"F593",X"F673",X"F754",X"F817",X"F8E1",X"F99D",X"FA23",X"FAA5",X"FB26",
		X"FBB7",X"FC6F",X"FD1F",X"FDD1",X"FE9F",X"FF67",X"0039",X"010A",X"01BB",X"027A",X"02FD",X"035E",X"0394",X"03AB",X"03AE",X"0397",
		X"035D",X"033B",X"034C",X"037D",X"03F0",X"0492",X"055D",X"064F",X"0779",X"08AE",X"09E7",X"0B10",X"0BE0",X"0C43",X"0C32",X"0BC4",
		X"0B31",X"0A8F",X"09A5",X"08BC",X"07D2",X"073D",X"06E8",X"06DD",X"0737",X"0773",X"07E0",X"0846",X"089D",X"08F0",X"0958",X"098E",
		X"098D",X"0947",X"08F8",X"08E5",X"0900",X"0938",X"098F",X"0A09",X"0A80",X"0B02",X"0BA1",X"0C2B",X"0C87",X"0CDD",X"0CA0",X"0C3B",
		X"0BB8",X"0B0A",X"0A73",X"09DF",X"0965",X"08E6",X"0859",X"0810",X"07EC",X"07D4",X"07CC",X"0777",X"0708",X"0656",X"0599",X"04B9",
		X"03B7",X"0293",X"0169",X"004A",X"FF3B",X"FE56",X"FDB5",X"FCFE",X"FC2E",X"FB77",X"FAAB",X"F9CB",X"F900",X"F838",X"F75F",X"F68D",
		X"F5A5",X"F4CF",X"F3DE",X"F319",X"F257",X"F1AA",X"F128",X"F0CE",X"F087",X"F04E",X"F03A",X"F016",X"F016",X"F00B",X"F01C",X"F03C",
		X"F053",X"F085",X"F0AE",X"F0BD",X"F0FA",X"F131",X"F174",X"F1CB",X"F21D",X"F274",X"F2C1",X"F335",X"F3A0",X"F423",X"F4B1",X"F545",
		X"F5DE",X"F662",X"F6E5",X"F771",X"F7D7",X"F840",X"F892",X"F902",X"F95F",X"F9C6",X"FA4D",X"FAFE",X"FBB1",X"FC69",X"FD4A",X"FE2E",
		X"FF32",X"001B",X"0103",X"01B2",X"0260",X"02F0",X"0373",X"03DE",X"0431",X"0464",X"0480",X"04AE",X"04F8",X"057D",X"0618",X"06C5",
		X"0795",X"083E",X"08F8",X"09B0",X"0A6C",X"0B3C",X"0BBE",X"0C33",X"0C5F",X"0C94",X"0CD4",X"0CFB",X"0D35",X"0D3D",X"0D53",X"0D72",
		X"0D6F",X"0D68",X"0D76",X"0D90",X"0D52",X"0D06",X"0C8D",X"0C09",X"0BC3",X"0B8D",X"0B67",X"0B23",X"0AD9",X"0ABE",X"0AA4",X"0A78",
		X"0A56",X"0A1C",X"09C9",X"0960",X"08F6",X"08AB",X"083B",X"07EA",X"0794",X"0749",X"0708",X"06C6",X"0692",X"066C",X"0644",X"0600",
		X"05A9",X"0528",X"049E",X"041A",X"03AF",X"031B",X"027B",X"01D3",X"012F",X"00A6",X"0032",X"FFAB",X"FEF8",X"FE4B",X"FD70",X"FCB1",
		X"FC15",X"FB80",X"FAE2",X"FA42",X"F9A8",X"F93A",X"F903",X"F8FE",X"F8F5",X"F8E8",X"F8B7",X"F86F",X"F83D",X"F7E2",X"F760",X"F6CE",
		X"F629",X"F579",X"F4DB",X"F448",X"F3E3",X"F394",X"F373",X"F34B",X"F347",X"F34F",X"F364",X"F38D",X"F3DE",X"F3F9",X"F405",X"F3EF",
		X"F406",X"F436",X"F457",X"F488",X"F4C4",X"F4F9",X"F559",X"F5CC",X"F650",X"F702",X"F7AA",X"F861",X"F8EF",X"F974",X"F9DF",X"FA3A",
		X"FA7D",X"FA9E",X"FAA7",X"FA93",X"FA7E",X"FA96",X"FABC",X"FAEF",X"FB3E",X"FBC9",X"FC5A",X"FCF7",X"FD89",X"FE15",X"FE87",X"FF0B",
		X"FF87",X"FFED",X"0054",X"00B2",X"00FF",X"0154",X"01C8",X"0234",X"02A0",X"0307",X"0361",X"03C4",X"0445",X"04D7",X"0567",X"05F1",
		X"0674",X"06F9",X"076B",X"07A6",X"07B6",X"07C3",X"079F",X"0769",X"0729",X"06CE",X"068E",X"069E",X"06E3",X"0729",X"0770",X"07C9",
		X"082B",X"086F",X"08A2",X"08A7",X"08AC",X"087F",X"0836",X"07E9",X"077C",X"0701",X"0691",X"064A",X"065A",X"0690",X"06BB",X"0709",
		X"074E",X"079E",X"07DA",X"0808",X"0821",X"07E9",X"07AB",X"0773",X"0748",X"0738",X"0715",X"0707",X"06E8",X"06F7",X"070C",X"0717",
		X"0719",X"06FF",X"06EA",X"06B5",X"0692",X"0672",X"064A",X"0623",X"05F7",X"05C1",X"0585",X"0533",X"04C1",X"044E",X"03DB",X"035F",
		X"02FA",X"0288",X"0206",X"0175",X"00CD",X"000A",X"FF04",X"FDF4",X"FCD1",X"FBB9",X"FAAF",X"F9A5",X"F8B3",X"F7EF",X"F761",X"F6DA",
		X"F66C",X"F5F6",X"F584",X"F530",X"F4F4",X"F4CE",X"F493",X"F43B",X"F410",X"F3CF",X"F3AF",X"F36D",X"F325",X"F2FD",X"F2E5",X"F2E9",
		X"F2C7",X"F2C5",X"F2EC",X"F32D",X"F378",X"F3E1",X"F447",X"F498",X"F51D",X"F5CA",X"F67D",X"F6FF",X"F78E",X"F7F2",X"F84E",X"F8B0",
		X"F90D",X"F94A",X"F956",X"F97C",X"F98D",X"F9C7",X"FA0C",X"FA4B",X"FAA8",X"FB09",X"FB75",X"FBEE",X"FC86",X"FCFB",X"FD54",X"FDB6",
		X"FE25",X"FE75",X"FEC0",X"FED5",X"FEC9",X"FE9E",X"FE58",X"FE22",X"FD9E",X"FD41",X"FCD3",X"FCA1",X"FCA5",X"FCB6",X"FD0B",X"FD6B",
		X"FE0F",X"FEE5",X"FFCD",X"00DF",X"01DF",X"02D3",X"03B6",X"04B3",X"05C2",X"06B3",X"079F",X"0888",X"0961",X"0A29",X"0B0F",X"0BD1",
		X"0CB2",X"0D68",X"0E2C",X"0EDF",X"0F69",X"0FE2",X"1047",X"1081",X"1086",X"1070",X"1055",X"102B",X"0FFB",X"1011",X"1051",X"1086",
		X"10BF",X"110E",X"114F",X"1182",X"119A",X"11AB",X"1182",X"113E",X"10D0",X"1054",X"0FCF",X"0F6B",X"0EEF",X"0E59",X"0DC7",X"0D3D",
		X"0CF4",X"0CBE",X"0C79",X"0C0C",X"0B5E",X"0A87",X"09C8",X"08E7",X"07BB",X"065B",X"04D9",X"0353",X"01D1",X"0083",X"FF2E",X"FDA7",
		X"FC59",X"FB2A",X"FA0D",X"F8FD",X"F828",X"F764",X"F68B",X"F5BF",X"F501",X"F467",X"F3B8",X"F31A",X"F28A",X"F210",X"F1B6",X"F143",
		X"F11F",X"F12E",X"F14C",X"F16E",X"F184",X"F1BB",X"F1B8",X"F1AD",X"F179",X"F152",X"F108",X"F096",X"F00F",X"EF80",X"EF28",X"EED7",
		X"EE7C",X"EE0B",X"EDA6",X"ED4E",X"ED11",X"ECE2",X"ECD5",X"ECC3",X"ECD4",X"ED23",X"ED93",X"EE0F",X"EE59",X"EEB3",X"EF19",X"EF75",
		X"EFD7",X"F028",X"F066",X"F0B0",X"F119",X"F195",X"F236",X"F2E0",X"F3D5",X"F4E2",X"F61D",X"F753",X"F875",X"F9A4",X"FABA",X"FBC1",
		X"FCC1",X"FDB6",X"FE9F",X"FF83",X"0056",X"014C",X"0245",X"034E",X"0462",X"0568",X"0677",X"0789",X"088A",X"0959",X"0A14",X"0ABD",
		X"0B64",X"0BE3",X"0C90",X"0D60",X"0E40",X"0F20",X"1039",X"1135",X"1242",X"1334",X"13FA",X"14AA",X"152D",X"1599",X"15C4",X"15DF",
		X"15B7",X"1594",X"1554",X"14FC",X"14C4",X"14A4",X"148B",X"1483",X"1467",X"1445",X"140F",X"13FC",X"13B7",X"1343",X"12B4",X"120F",
		X"1152",X"1089",X"0FB6",X"0EF5",X"0E46",X"0D6B",X"0CBC",X"0C10",X"0B5E",X"0AC7",X"0A3F",X"09B3",X"0900",X"0875",X"07F2",X"0761",
		X"06C5",X"0626",X"0556",X"0493",X"03C3",X"02D8",X"0207",X"012E",X"0059",X"FF52",X"FE3F",X"FD46",X"FC69",X"FBC8",X"FB11",X"FA58",
		X"F993",X"F8D1",X"F812",X"F785",X"F6FA",X"F626",X"F540",X"F459",X"F39A",X"F2D3",X"F21B",X"F159",X"F099",X"EFBE",X"EF23",X"EEAD",
		X"EE2F",X"ED9F",X"ED22",X"ECED",X"ECBB",X"EC68",X"EC1A",X"EBD8",X"EBB5",X"EB99",X"EB70",X"EB60",X"EB4C",X"EB57",X"EB78",X"EB9A",
		X"EBF7",X"EC59",X"ECBD",X"ED2A",X"ED85",X"EE14",X"EE96",X"EF06",X"EF98",X"F006",X"F07E",X"F119",X"F1B5",X"F245",X"F2C9",X"F35F",
		X"F3F3",X"F4B0",X"F583",X"F65F",X"F73E",X"F82E",X"F94D",X"FA57",X"FB5A",X"FC64",X"FD86",X"FE7B",X"FF31",X"FFE3",X"00AB",X"0169",
		X"021C",X"02D5",X"0395",X"042F",X"04E8",X"05EF",X"06F4",X"07F8",X"08F4",X"09FB",X"0ADD",X"0B8E",X"0C2B",X"0C9D",X"0CDB",X"0CEA",
		X"0CBE",X"0C9F",X"0C8B",X"0C7F",X"0C89",X"0CCA",X"0D5E",X"0E2F",X"0F20",X"1014",X"1107",X"11F4",X"12CE",X"1363",X"13B7",X"13DA",
		X"13F1",X"13CF",X"1388",X"1361",X"1344",X"1344",X"135C",X"137C",X"1387",X"1383",X"1382",X"135D",X"12E7",X"123A",X"1174",X"10A3",
		X"0FA0",X"0EAB",X"0DE7",X"0D1E",X"0C71",X"0BFC",X"0B8D",X"0B54",X"0B12",X"0AC8",X"0A3D",X"09A0",X"0914",X"0850",X"0721",X"05FD",
		X"04C1",X"039D",X"0295",X"0195",X"00C0",X"FFF8",X"FF56",X"FEBF",X"FE45",X"FDBF",X"FD4D",X"FCEE",X"FC72",X"FBB4",X"FAF6",X"FA28",
		X"F959",X"F88A",X"F7B2",X"F6D4",X"F60A",X"F566",X"F4D3",X"F453",X"F3FF",X"F392",X"F351",X"F321",X"F319",X"F316",X"F31D",X"F2FA",
		X"F2C0",X"F2A0",X"F271",X"F24C",X"F223",X"F202",X"F1BF",X"F169",X"F121",X"F0F3",X"F0B7",X"F05C",X"EFD3",X"EF6F",X"EF17",X"EEBB",
		X"EE6D",X"EE44",X"EE1F",X"EDF5",X"EDB7",X"ED90",X"ED6F",X"ED51",X"ED6C",X"ED9C",X"EDDD",X"EE1F",X"EE66",X"EED3",X"EF51",X"EFCA",
		X"F071",X"F132",X"F205",X"F2E0",X"F3D7",X"F4EE",X"F5F5",X"F6F5",X"F7DF",X"F8B6",X"F97D",X"FA61",X"FB1C",X"FBE6",X"FCBE",X"FD93",
		X"FE88",X"FF79",X"007E",X"0187",X"0270",X"0360",X"0456",X"052C",X"05FA",X"06A7",X"073C",X"07BA",X"0813",X"089C",X"0940",X"09A8",
		X"0A16",X"0A8B",X"0B07",X"0B9E",X"0C22",X"0CA8",X"0D2C",X"0D8A",X"0DF0",X"0E38",X"0E72",X"0EB0",X"0EDD",X"0EFC",X"0F08",X"0F08",
		X"0F29",X"0F1B",X"0F1D",X"0F4A",X"0F8C",X"0FC5",X"0FF6",X"1025",X"1046",X"104F",X"1032",X"100A",X"0F92",X"0EED",X"0E63",X"0DDE",
		X"0D6E",X"0D01",X"0CB6",X"0C8E",X"0C93",X"0CBE",X"0D16",X"0D89",X"0DCA",X"0DF0",X"0DC8",X"0D69",X"0CF6",X"0C70",X"0BA4",X"0AAA",
		X"0996",X"0874",X"076A",X"0676",X"05A4",X"0502",X"0459",X"03DB",X"033B",X"02AC",X"0212",X"017C",X"0100",X"0078",X"FFD1",X"FF29",
		X"FE89",X"FDF6",X"FDA9",X"FD59",X"FD09",X"FCA1",X"FC46",X"FC04",X"FBF8",X"FBEB",X"FBB1",X"FB62",X"FB01",X"FA9E",X"FA4F",X"F9D8",
		X"F92D",X"F87E",X"F7BF",X"F6F4",X"F624",X"F575",X"F4F1",X"F467",X"F3E5",X"F38E",X"F35A",X"F34E",X"F353",X"F37D",X"F382",X"F366",
		X"F355",X"F326",X"F2EA",X"F2A9",X"F23C",X"F1B0",X"F111",X"F07B",X"F015",X"EFDF",X"EFEC",X"F005",X"F033",X"F075",X"F0E3",X"F15F",
		X"F1EA",X"F25B",X"F2AB",X"F2D4",X"F29C",X"F279",X"F270",X"F26A",X"F264",X"F261",X"F291",X"F2CA",X"F337",X"F3C0",X"F466",X"F51D",
		X"F5F2",X"F6C6",X"F7C5",X"F8AE",X"F9A8",X"FA71",X"FB18",X"FBB4",X"FC51",X"FCEA",X"FD7F",X"FE24",X"FED1",X"FF7F",X"0031",X"00E9",
		X"0172",X"021E",X"02A5",X"0335",X"03A0",X"0408",X"0463",X"04AB",X"0503",X"0571",X"05FB",X"0682",X"0733",X"0809",X"08F9",X"09DA",
		X"0A91",X"0B55",X"0BE9",X"0C5A",X"0CA2",X"0CB9",X"0C7C",X"0C2D",X"0BA1",X"0AFA",X"0A7E",X"0A01",X"09DC",X"09E0",X"09F6",X"0A39",
		X"0AB7",X"0B62",X"0C2A",X"0D07",X"0DDF",X"0E82",X"0F00",X"0F71",X"0FB5",X"0FE6",X"1001",X"0FEE",X"0FC8",X"0FA0",X"0F87",X"0F7F",
		X"0F97",X"0F99",X"0FB7",X"0FDB",X"1008",X"1032",X"1038",X"102A",X"0FD3",X"0F50",X"0EAB",X"0DE7",X"0D37",X"0C75",X"0BB3",X"0B2F",
		X"0ABA",X"0A3C",X"09C1",X"0979",X"0921",X"08B4",X"0865",X"07F3",X"075E",X"069D",X"05CF",X"0506",X"0401",X"030F",X"0225",X"014D",
		X"007F",X"FFAA",X"FED1",X"FDEC",X"FCC4",X"FB94",X"FA5C",X"F912",X"F7D1",X"F684",X"F558",X"F430",X"F300",X"F1F1",X"F0E5",X"F00C",
		X"EF21",X"EE19",X"ED3D",X"EC75",X"EBBF",X"EB3E",X"EAD7",X"EA7B",X"EA33",X"EA07",X"E9EF",X"E9F4",X"EA21",X"EA5B",X"EAB1",X"EAE7",
		X"EB43",X"EBCB",X"EC57",X"ECB4",X"ED25",X"ED97",X"EE0E",X"EE61",X"EEBB",X"EF11",X"EF3A",X"EF5B",X"EF7B",X"EFA6",X"EFB7",X"EFB8",
		X"EFC4",X"EFCB",X"F002",X"F05D",X"F0D4",X"F183",X"F243",X"F30D",X"F3F3",X"F4D8",X"F5C3",X"F6BD",X"F7BB",X"F8BC",X"F9A3",X"FAAF",
		X"FBA1",X"FC6C",X"FD3C",X"FE41",X"FF48",X"004A",X"013F",X"0268",X"03A5",X"04D5",X"0611",X"0754",X"0877",X"095B",X"0A6B",X"0B65",
		X"0C30",X"0CB7",X"0D2B",X"0D8E",X"0DE2",X"0E1D",X"0E54",X"0E73",X"0EA4",X"0EF7",X"0F46",X"0FB7",X"104B",X"10E4",X"1186",X"1240",
		X"12F5",X"13A6",X"1441",X"14E3",X"156A",X"15FE",X"1679",X"16E4",X"16F9",X"1702",X"16FD",X"16E7",X"16C0",X"1680",X"164A",X"15F8",
		X"15A9",X"157C",X"155B",X"1508",X"148F",X"13F9",X"1343",X"128C",X"11A0",X"10B1",X"0FA2",X"0E6F",X"0D2F",X"0BF0",X"0AC4",X"09B5",
		X"08E9",X"083C",X"078D",X"06E4",X"0636",X"0569",X"0483",X"0391",X"026B",X"0147",X"0002",X"FEA0",X"FD5B",X"FC30",X"FB38",X"FA47",
		X"F98A",X"F8DE",X"F865",X"F7DC",X"F764",X"F6B1",X"F5EC",X"F50B",X"F3FA",X"F2F0",X"F1D6",X"F0BB",X"EFA5",X"EE94",X"ED95",X"ECC4",
		X"EC14",X"EB9D",X"EB3C",X"EABF",X"EA6B",X"EA21",X"E9DB",X"E97C",X"E923",X"E8E8",X"E8B6",X"E898",X"E873",X"E85C",X"E86C",X"E8A3",
		X"E8D3",X"E936",X"E96D",X"E9AC",X"E9F5",X"EA2D",X"EA5E",X"EA69",X"EA9E",X"EA9D",X"EACC",X"EB11",X"EB47",X"EB9B",X"EC29",X"ECF3",
		X"EDEE",X"EF45",X"F0C0",X"F267",X"F409",X"F5C8",X"F78C",X"F95C",X"FB1E",X"FCB7",X"FE1A",X"FF53",X"0088",X"0199",X"02B1",X"03A5",
		X"046A",X"0538",X"0605",X"06F8",X"07F0",X"08DD",X"09C4",X"0AA3",X"0BBF",X"0CDA",X"0E15",X"0F48",X"1082",X"11BA",X"12E0",X"13F2",
		X"14F0",X"15EC",X"1694",X"171F",X"17A2",X"1820",X"1891",X"1904",X"1960",X"19B0",X"19E6",X"19F6",X"1A10",X"1A17",X"19E4",X"198D",
		X"190E",X"1865",X"1796",X"16AF",X"15CB",X"14FA",X"142A",X"135A",X"1295",X"121A",X"11A0",X"1141",X"10CE",X"1025",X"0F6F",X"0EC0",
		X"0E28",X"0D4F",X"0C63",X"0B5B",X"0A23",X"090D",X"0828",X"0723",X"0607",X"04FE",X"03F4",X"02D3",X"01A1",X"0070",X"FF48",X"FDE3",
		X"FCA7",X"FB6C",X"FA45",X"F95E",X"F896",X"F806",X"F77A",X"F6E8",X"F6AD",X"F66A",X"F647",X"F63A",X"F62A",X"F60B",X"F5D8",X"F578",
		X"F509",X"F4A2",X"F418",X"F3A3",X"F319",X"F28E",X"F20B",X"F1B3",X"F15B",X"F11A",X"F0CC",X"F0A8",X"F094",X"F095",X"F09B",X"F06B",
		X"F06E",X"F058",X"F040",X"F01E",X"EFFD",X"EFE6",X"EFEA",X"EFD9",X"EFE4",X"F00B",X"F048",X"F09B",X"F11C",X"F1B2",X"F21F",X"F28A",
		X"F2CE",X"F31A",X"F33F",X"F351",X"F337",X"F300",X"F2D5",X"F283",X"F245",X"F202",X"F1F7",X"F222",X"F253",X"F291",X"F2F6",X"F397",
		X"F437",X"F4E5",X"F5CD",X"F6AB",X"F76B",X"F83B",X"F8F9",X"F9C9",X"FA92",X"FB65",X"FC32",X"FCFA",X"FDCC",X"FE79",X"FF04",X"FFC2",
		X"0083",X"0106",X"017C",X"01E5",X"027F",X"0329",X"0410",X"050E",X"05F4",X"06CE",X"07B9",X"08CD",X"09CF",X"0AD0",X"0B98",X"0C54",
		X"0CFF",X"0DC8",X"0EA1",X"0F7D",X"106D",X"1172",X"126B",X"134F",X"1445",X"150F",X"159E",X"15FA",X"15F8",X"15DF",X"15C6",X"1597",
		X"1562",X"1516",X"14D4",X"149D",X"148A",X"149B",X"14CD",X"1507",X"151A",X"152D",X"1541",X"1528",X"14ED",X"14A0",X"1438",X"1394",
		X"1314",X"1276",X"11CF",X"112B",X"1090",X"0FD9",X"0F16",X"0E4A",X"0D5E",X"0C36",X"0ABE",X"093E",X"0795",X"05F9",X"0459",X"02D6",
		X"016F",X"0022",X"FF0B",X"FE0B",X"FD32",X"FC6E",X"FBE4",X"FB4B",X"FA8D",X"F998",X"F891",X"F77E",X"F647",X"F502",X"F3AD",X"F272",
		X"F15A",X"F07A",X"EFCB",X"EF42",X"EEBC",X"EE64",X"EE4A",X"EE39",X"EE3A",X"EE3B",X"EE19",X"EDF7",X"EDDE",X"ED92",X"ED25",X"ECD5",
		X"EC99",X"EC6C",X"EC70",X"ECAE",X"ED02",X"ED50",X"EDA9",X"EE24",X"EEB2",X"EF45",X"EFB7",X"F013",X"F05D",X"F0AC",X"F0E8",X"F116",
		X"F16C",X"F1DB",X"F251",X"F2C9",X"F33E",X"F3C3",X"F465",X"F510",X"F5B2",X"F614",X"F648",X"F69A",X"F6F9",X"F779",X"F7FD",X"F852",
		X"F8B9",X"F914",X"F973",X"FA08",X"FA76",X"FAEC",X"FB33",X"FB73",X"FBE4",X"FC3D",X"FCC9",X"FD76",X"FE29",X"FF05",X"0004",X"0105",
		X"021C",X"033B",X"0456",X"0548",X"060B",X"06A6",X"0723",X"07A5",X"0839",X"08DB",X"0959",X"09EA",X"0A93",X"0B4E",X"0C21",X"0CF5",
		X"0DC0",X"0E9E",X"0F5B",X"1017",X"10E6",X"11A1",X"1240",X"12D6",X"1349",X"1385",X"13AC",X"13FE",X"1436",X"1447",X"144A",X"1406",
		X"13B8",X"1368",X"1338",X"12F6",X"12BC",X"1280",X"124F",X"122E",X"1208",X"1217",X"1233",X"1235",X"1200",X"11CB",X"117D",X"10D7",
		X"0FFE",X"0F11",X"0E13",X"0CFE",X"0BDB",X"0A9C",X"094E",X"080E",X"06EF",X"05C3",X"0474",X"030E",X"01AB",X"0056",X"FF09",X"FDD8",
		X"FCBB",X"FBA0",X"FA8D",X"F9C3",X"F924",X"F882",X"F7FB",X"F774",X"F6DD",X"F64D",X"F5E6",X"F568",X"F4CE",X"F42E",X"F374",X"F2DC",
		X"F241",X"F1A8",X"F142",X"F0DC",X"F083",X"F050",X"F063",X"F0A4",X"F0D4",X"F102",X"F114",X"F0FA",X"F0D9",X"F09D",X"F027",X"EFB7",
		X"EF3A",X"EEDD",X"EEA5",X"EE93",X"EEBE",X"EEE8",X"EF3F",X"EFBA",X"F025",X"F087",X"F0BF",X"F112",X"F185",X"F1D3",X"F225",X"F26F",
		X"F2A2",X"F2E9",X"F362",X"F3F1",X"F470",X"F4F0",X"F576",X"F5FD",X"F664",X"F6AA",X"F6C3",X"F6AD",X"F68C",X"F685",X"F6CB",X"F700",
		X"F781",X"F831",X"F90E",X"FA1A",X"FB46",X"FC8C",X"FDF5",X"FF4B",X"00AD",X"0224",X"0388",X"04D6",X"05D7",X"06D1",X"07A6",X"0869",
		X"091A",X"09C1",X"0A3A",X"0AE1",X"0B82",X"0C0C",X"0C9B",X"0D16",X"0D71",X"0DD6",X"0E48",X"0EB2",X"0F28",X"0F7F",X"1002",X"1060",
		X"10F6",X"1197",X"1211",X"1294",X"12F6",X"134E",X"1382",X"13A5",X"13AE",X"13C5",X"13A6",X"1369",X"1311",X"129E",X"1200",X"116C",
		X"10D2",X"1039",X"0F9B",X"0F07",X"0E88",X"0E0B",X"0D7C",X"0CF2",X"0C75",X"0BCA",X"0B18",X"0A3F",X"0970",X"08BB",X"07F3",X"0740",
		X"06A3",X"05D6",X"04F0",X"03FC",X"0314",X"0217",X"012F",X"005B",X"FFA1",X"FEFD",X"FE79",X"FE15",X"FDC8",X"FD73",X"FD07",X"FC9A",
		X"FC02",X"FB4B",X"FAA3",X"F9D1",X"F900",X"F855",X"F798",X"F6E0",X"F62F",X"F5CB",X"F574",X"F54F",X"F533",X"F517",X"F4D8",X"F493",
		X"F445",X"F3CC",X"F35A",X"F2F3",X"F2A0",X"F24E",X"F203",X"F1C6",X"F1B4",X"F19D",X"F1C3",X"F1CD",X"F1C3",X"F19C",X"F162",X"F12C",
		X"F0F0",X"F0C0",X"F086",X"F06F",X"F083",X"F0ED",X"F175",X"F200",X"F2A5",X"F360",X"F41D",X"F4D4",X"F58D",X"F623",X"F6B1",X"F726",
		X"F7B2",X"F81A",X"F869",X"F8D1",X"F924",X"F95A",X"F991",X"F9CD",X"FA19",X"FA66",X"FADE",X"FB56",X"FBCB",X"FC44",X"FCA2",X"FD2E",
		X"FDB5",X"FE3D",X"FECB",X"FF45",X"FF9D",X"0006",X"00A4",X"0152",X"020C",X"02AD",X"034F",X"0403",X"04CE",X"0597",X"0663",X"073E",
		X"07EA",X"08AC",X"0973",X"0A2C",X"0AE3",X"0B89",X"0C4B",X"0D00",X"0DA8",X"0E1D",X"0E89",X"0EF6",X"0F54",X"0F90",X"0FD7",X"1014",
		X"104A",X"10B2",X"10FD",X"1136",X"1144",X"117A",X"11B6",X"1210",X"126C",X"127A",X"126A",X"124E",X"1230",X"1209",X"1195",X"1116",
		X"10A8",X"100D",X"0F81",X"0EEC",X"0E52",X"0DA0",X"0CB9",X"0BC7",X"0AA9",X"097A",X"084E",X"06FC",X"05D3",X"04DF",X"03EE",X"02DC",
		X"01BB",X"00BA",X"FFCB",X"FEFB",X"FE0E",X"FD00",X"FBB2",X"FA51",X"F914",X"F7F1",X"F6CC",X"F5B6",X"F4B4",X"F3B7",X"F302",X"F291",
		X"F21F",X"F1A6",X"F12F",X"F0CA",X"F056",X"EFD5",X"EF62",X"EEE9",X"EE71",X"EE0A",X"EDAF",X"ED62",X"ED72",X"EDBA",X"EE2D",X"EECB",
		X"EF69",X"F00D",X"F08F",X"F133",X"F1DB",X"F276",X"F2DF",X"F31A",X"F33B",X"F365",X"F39D",X"F411",X"F486",X"F50B",X"F569",X"F609",
		X"F6E3",X"F7CC",X"F8C5",X"F99E",X"FA69",X"FB09",X"FBB7",X"FC4A",X"FCC3",X"FD21",X"FD82",X"FDDD",X"FE29",X"FE81",X"FF05",X"FFAA",
		X"006B",X"0134",X"0203",X"02BC",X"037B",X"0455",X"051D",X"05CF",X"065F",X"06CB",X"072E",X"077D",X"07D7",X"0827",X"0863",X"08A0",
		X"08CC",X"08ED",X"0902",X"090D",X"08F8",X"08B9",X"087F",X"083A",X"07EB",X"07B0",X"0787",X"0767",X"0762",X"077D",X"07B2",X"0813",
		X"0887",X"08F3",X"0947",X"096E",X"096F",X"0980",X"095B",X"0929",X"08E4",X"0898",X"0854",X"07EA",X"0791",X"0761",X"0731",X"06EB",
		X"06B0",X"067A",X"0660",X"0657",X"066B",X"0675",X"066F",X"065D",X"0658",X"0654",X"0637",X"060C",X"05CA",X"057C",X"051C",X"04BB",
		X"045E",X"0401",X"03E3",X"039E",X"035B",X"030B",X"02CE",X"028E",X"0218",X"01B4",X"0135",X"00B0",X"0005",X"FF6B",X"FEDF",X"FE4F",
		X"FDC8",X"FD5B",X"FCEA",X"FC86",X"FC3A",X"FBEA",X"FB81",X"FAF2",X"FA64",X"F9BF",X"F8ED",X"F84E",X"F7B8",X"F726",X"F6BC",X"F659",
		X"F636",X"F61A",X"F616",X"F628",X"F62C",X"F646",X"F67D",X"F6A3",X"F6AD",X"F697",X"F675",X"F64B",X"F631",X"F60C",X"F5F6",X"F624",
		X"F62B",X"F64E",X"F6B1",X"F711",X"F763",X"F7D0",X"F82D",X"F8A4",X"F932",X"F9C2",X"FA4F",X"FAE2",X"FB70",X"FC28",X"FCCE",X"FD53",
		X"FDD1",X"FE33",X"FEA1",X"FEC1",X"FEE7",X"FEE3",X"FEAA",X"FE73",X"FE7B",X"FE8E",X"FE89",X"FE95",X"FEAA",X"FEE6",X"FF1F",X"FF55",
		X"FF68",X"FF67",X"FF2E",X"FEFA",X"FEBA",X"FE9E",X"FEA8",X"FEC4",X"FF35",X"FFB2",X"0066",X"0141",X"0224",X"02F6",X"03A9",X"043C",
		X"04B2",X"04E9",X"0512",X"0523",X"04FD",X"04E2",X"048D",X"043F",X"041B",X"041B",X"0493",X"052A",X"05CF",X"0656",X"06EE",X"079F",
		X"0859",X"0903",X"0966",X"098A",X"0957",X"091B",X"08C2",X"0884",X"0830",X"07B9",X"0778",X"0750",X"075E",X"0778",X"079D",X"0795",
		X"076D",X"0773",X"0755",X"074D",X"0727",X"070B",X"06BE",X"0672",X"061D",X"05E2",X"05C8",X"05B7",X"05A0",X"054C",X"04D9",X"045D",
		X"03FD",X"0356",X"02A2",X"01EB",X"0158",X"00D9",X"007F",X"003C",X"0027",X"002E",X"004E",X"0052",X"005C",X"0073",X"006A",X"0070",
		X"003F",X"FFEE",X"FF68",X"FEE1",X"FE8D",X"FE36",X"FDE2",X"FDA6",X"FD77",X"FD40",X"FD11",X"FD09",X"FD22",X"FCE6",X"FC74",X"FBF0",
		X"FB50",X"FAC6",X"FA5E",X"F9F6",X"F989",X"F91F",X"F8AB",X"F87B",X"F83C",X"F808",X"F7E2",X"F7AE",X"F77E",X"F75F",X"F774",X"F76D",
		X"F734",X"F6DE",X"F6A0",X"F64C",X"F612",X"F5E3",X"F5AE",X"F57B",X"F567",X"F589",X"F5BC",X"F606",X"F657",X"F6CF",X"F72E",X"F7A2",
		X"F836",X"F8BF",X"F93C",X"F976",X"F9CA",X"FA19",X"FA54",X"FAC2",X"FB3F",X"FBC1",X"FC69",X"FD23",X"FDCF",X"FE84",X"FF47",X"0011",
		X"00AE",X"0127",X"019C",X"01FA",X"023C",X"02BE",X"0338",X"03A4",X"0422",X"0494",X"0520",X"05B9",X"0669",X"070F",X"0791",X"07EB",
		X"083A",X"0888",X"0892",X"0870",X"0831",X"07E3",X"0794",X"0754",X"0743",X"0714",X"0716",X"0752",X"0786",X"07DA",X"0834",X"0883",
		X"08B2",X"0899",X"089D",X"086C",X"07FB",X"0772",X"06D8",X"063A",X"0588",X"0501",X"04A9",X"042F",X"03CC",X"03A1",X"0392",X"03AF",
		X"03CB",X"03CB",X"03B8",X"03B8",X"03C8",X"03C3",X"03B7",X"03C1",X"03A5",X"0398",X"0369",X"0335",X"02EF",X"02AD",X"0251",X"01E8",
		X"0188",X"00D9",X"004F",X"FFAA",X"FF00",X"FE5E",X"FDC2",X"FD15",X"FC94",X"FC18",X"FBB5",X"FB5F",X"FAF3",X"FA8E",X"FA58",X"FA35",
		X"FA08",X"F9F5",X"F9CE",X"F99C",X"F983",X"F96C",X"F95F",X"F967",X"F970",X"F978",X"F950",X"F95E",X"F992",X"F9C0",X"F9E6",X"F9F9",
		X"FA11",X"FA28",X"FA3C",X"FA5F",X"FA77",X"FA8F",X"FACD",X"FAEB",X"FAFA",X"FB28",X"FB55",X"FB80",X"FBA7",X"FBD8",X"FBE4",X"FC13",
		X"FC63",X"FCB5",X"FD2C",X"FD81",X"FDC6",X"FE17",X"FE77",X"FF02",X"FF65",X"FFCE",X"0008",X"0047",X"00B6",X"0123",X"0187",X"01D6",
		X"0218",X"0273",X"02E9",X"0340",X"0384",X"03B3",X"03C6",X"03F9",X"0419",X"0422",X"042B",X"044F",X"0465",X"0495",X"04BE",X"04DC",
		X"051C",X"0572",X"05D5",X"0618",X"0653",X"0645",X"0649",X"063A",X"05EA",X"059F",X"0552",X"04C7",X"043A",X"03AD",X"0354",X"02F4",
		X"02AD",X"0277",X"0251",X"0254",X"0269",X"028C",X"02A4",X"02AF",X"02C3",X"02B5",X"0296",X"0256",X"020A",X"01BC",X"0153",X"0117",
		X"00CE",X"0097",X"007F",X"007C",X"0076",X"007F",X"0087",X"00AC",X"00AF",X"0072",X"002C",X"FFBC",X"FF43",X"FED3",X"FE2E",X"FD85",
		X"FCE6",X"FC50",X"FC00",X"FB7C",X"FB2D",X"FAEE",X"FAF3",X"FB17",X"FB34",X"FB6F",X"FB8F",X"FBCF",X"FC16",X"FC52",X"FC6F",X"FC84",
		X"FC8C",X"FCBC",X"FCEE",X"FD35",X"FD59",X"FD51",X"FD57",X"FD2D",X"FD1B",X"FD07",X"FCAD",X"FC48",X"FBFE",X"FB9C",X"FB6E",X"FB40",
		X"FAFF",X"FACC",X"FAA3",X"FA8B",X"FA95",X"FABA",X"FB10",X"FB5A",X"FBA4",X"FC36",X"FCC6",X"FD5F",X"FDDA",X"FE60",X"FEDF",X"FF80",
		X"FFFF",X"0087",X"00CE",X"010F",X"0176",X"01DC",X"024D",X"02B0",X"030F",X"0364",X"03CB",X"043E",X"04A2",X"04C5",X"04CF",X"04E2",
		X"04BF",X"04B8",X"049D",X"0453",X"0410",X"03E3",X"03BE",X"03C2",X"03CF",X"039E",X"037E",X"033B",X"02EC",X"02A9",X"023F",X"01CE",
		X"0153",X"00F0",X"00A5",X"008D",X"0081",X"0099",X"00BD",X"00E2",X"0112",X"0121",X"0157",X"017F",X"01BC",X"01BC",X"01A3",X"0199",
		X"018A",X"017D",X"0162",X"013C",X"0128",X"0114",X"012D",X"0174",X"01AA",X"01CE",X"01E8",X"01FF",X"0226",X"0219",X"0233",X"01F8",
		X"01A3",X"0171",X"014B",X"0120",X"010C",X"012F",X"015F",X"018B",X"01D6",X"0255",X"02B4",X"0307",X"0360",X"0380",X"0377",X"036E",
		X"034A",X"0306",X"0294",X"0211",X"019E",X"0143",X"00E3",X"00C8",X"00A7",X"0069",X"003B",X"0004",X"FFA9",X"FF42",X"FED5",X"FE47",
		X"FD89",X"FCE9",X"FC50",X"FBD6",X"FB7B",X"FB3B",X"FAF7",X"FAB1",X"FA9B",X"FA85",X"FA68",X"FA53",X"FA43",X"FA2B",X"FA13",X"FA08",
		X"F9FE",X"FA2B",X"FA72",X"FAC6",X"FB0B",X"FB2E",X"FB75",X"FBA2",X"FBBA",X"FBAA",X"FB75",X"FB0C",X"FA92",X"F9E6",X"F951",X"F8CE",
		X"F886",X"F83C",X"F81C",X"F82E",X"F889",X"F90B",X"F9BB",X"FA6C",X"FAF9",X"FB84",X"FC2F",X"FCBC",X"FD40",X"FDD5",X"FE45",X"FE90",
		X"FEF1",X"FF62",X"FFBD",X"002C",X"00B2",X"0142",X"01C0",X"023B",X"0284",X"02E9",X"0334",X"0369",X"0375",X"0372",X"034F",X"033C",
		X"0373",X"03A1",X"040E",X"0467",X"04ED",X"055B",X"05F1",X"06B3",X"072A",X"079C",X"07DA",X"07FF",X"07E7",X"07F0",X"07ED",X"07D3",
		X"07B0",X"07B1",X"07EF",X"0811",X"084F",X"087E",X"08B3",X"08D8",X"08D5",X"08D8",X"08B1",X"0865",X"07E6",X"0771",X"06E6",X"065A",
		X"05CA",X"054C",X"04D0",X"0497",X"0464",X"042B",X"03EE",X"03A4",X"0369",X"0330",X"0305",X"02C7",X"0253",X"0201",X"01B7",X"017B",
		X"0180",X"0144",X"00EF",X"008F",X"002D",X"FFED",X"FF9D",X"FF3E",X"FEBD",X"FE32",X"FDAB",X"FD53",X"FD08",X"FCA8",X"FC63",X"FC1B",
		X"FBDE",X"FB87",X"FB78",X"FB64",X"FB3E",X"FB1F",X"FAF0",X"FABC",X"FA96",X"FA8D",X"FA8B",X"FA5F",X"FA35",X"FA07",X"F9C2",X"F9AE",
		X"F9C0",X"F9BB",X"F983",X"F96D",X"F945",X"F945",X"F943",X"F941",X"F93A",X"F91C",X"F90E",X"F923",X"F93A",X"F94A",X"F97E",X"F984",
		X"F9B3",X"F9D2",X"FA19",X"FA67",X"FA8E",X"FAD3",X"FAF7",X"FB29",X"FB43",X"FB52",X"FB6A",X"FB61",X"FB79",X"FB72",X"FB88",X"FB9C",
		X"FBB6",X"FBD9",X"FBE8",X"FBC7",X"FB97",X"FB78",X"FB42",X"FB34",X"FB5B",X"FBBD",X"FC2C",X"FCCB",X"FD6D",X"FE47",X"FF25",X"FFFD",
		X"00B5",X"011B",X"0168",X"01D4",X"0250",X"02A9",X"035C",X"0410",X"04E2",X"05D3",X"06E4",X"0807",X"08FF",X"09D5",X"0A75",X"0AFE",
		X"0B28",X"0B39",X"0B3F",X"0B4D",X"0B46",X"0B42",X"0B60",X"0B73",X"0B94",X"0BDF",X"0C37",X"0C42",X"0C28",X"0C1F",X"0BF5",X"0BB6",
		X"0B75",X"0AF7",X"0A63",X"09D7",X"0962",X"0924",X"08F8",X"08C9",X"08A4",X"0888",X"0854",X"0826",X"07F2",X"0797",X"0701",X"063E",
		X"0554",X"043F",X"0343",X"022D",X"00EC",X"FFB3",X"FEAD",X"FD9E",X"FC8F",X"FB8C",X"FAD8",X"FA0E",X"F960",X"F8B0",X"F808",X"F767",
		X"F6D5",X"F666",X"F5D2",X"F564",X"F4F4",X"F4AC",X"F472",X"F439",X"F418",X"F3E8",X"F3AA",X"F380",X"F343",X"F330",X"F327",X"F311",
		X"F2F0",X"F2DE",X"F302",X"F320",X"F344",X"F383",X"F3C0",X"F411",X"F453",X"F49E",X"F4B5",X"F4C9",X"F4DB",X"F4C9",X"F4AB",X"F486",
		X"F494",X"F4A4",X"F4DF",X"F52B",X"F5B7",X"F66D",X"F70C",X"F800",X"F8E3",X"F9A7",X"FAAE",X"FB83",X"FC18",X"FCC5",X"FD78",X"FE42",
		X"FEF0",X"FFB6",X"009E",X"016A",X"025C",X"0362",X"044C",X"04F5",X"057F",X"062C",X"06B0",X"06F3",X"0760",X"07D5",X"0852",X"08E2",
		X"0974",X"0A01",X"0A90",X"0B37",X"0BE9",X"0C8B",X"0D0A",X"0D6A",X"0DBD",X"0DEE",X"0E23",X"0E5B",X"0E7D",X"0EB2",X"0EF9",X"0F56",
		X"0F9F",X"0FE7",X"101F",X"105D",X"1082",X"1076",X"1064",X"1040",X"100B",X"0FCB",X"0F88",X"0F45",X"0F15",X"0EB2",X"0E46",X"0DAC",
		X"0D1B",X"0C55",X"0B60",X"0A6D",X"095F",X"083E",X"071E",X"062F",X"054A",X"045D",X"039A",X"0313",X"02B9",X"027D",X"0232",X"01C9",
		X"0183",X"012C",X"009C",X"000F",X"FF60",X"FEA3",X"FE05",X"FD70",X"FCF2",X"FC85",X"FC05",X"FB9B",X"FB42",X"FAB7",X"FA0E",X"F940",
		X"F862",X"F74B",X"F63C",X"F52B",X"F41E",X"F35B",X"F292",X"F202",X"F187",X"F13F",X"F10D",X"F0FD",X"F0CA",X"F0AD",X"F081",X"F037",
		X"EFFD",X"EFBF",X"EF98",X"EF67",X"EF53",X"EF0D",X"EEDF",X"EED5",X"EEE0",X"EF1C",X"EF48",X"EF94",X"EFC8",X"EFF9",X"F036",X"F06F",
		X"F0AB",X"F0B5",X"F0CA",X"F102",X"F127",X"F18A",X"F201",X"F2A0",X"F341",X"F3F1",X"F4A4",X"F55B",X"F628",X"F714",X"F800",X"F8E0",
		X"F9CC",X"FABB",X"FBDC",X"FD2E",X"FE85",X"FFC8",X"00ED",X"01D3",X"02E6",X"0400",X"0523",X"064D",X"0756",X"085C",X"0964",X"0A59",
		X"0B5C",X"0C3A",X"0CEB",X"0D64",X"0DB2",X"0E0F",X"0E89",X"0F01",X"0F6C",X"0FE0",X"1038",X"109B",X"1138",X"11CE",X"1275",X"1314",
		X"139F",X"1421",X"149B",X"151A",X"1580",X"15D2",X"15FB",X"1601",X"1616",X"1612",X"1632",X"1636",X"1620",X"1616",X"15C4",X"1583",
		X"153A",X"14E4",X"1476",X"13D1",X"12DE",X"11E3",X"10C9",X"0F92",X"0E60",X"0CF6",X"0B6A",X"09BF",X"0836",X"06C0",X"055F",X"0405",
		X"02B9",X"016F",X"0029",X"FF15",X"FE20",X"FD2E",X"FC0C",X"FB07",X"FA04",X"F912",X"F823",X"F731",X"F65E",X"F583",X"F4CB",X"F3F7",
		X"F320",X"F256",X"F183",X"F0A3",X"EFB9",X"EEC9",X"EDD1",X"ECDC",X"EBE6",X"EB06",X"EA25",X"E948",X"E862",X"E78B",X"E6FD",X"E6AA",
		X"E67E",X"E65C",X"E674",X"E6D9",X"E76A",X"E84A",X"E931",X"EA2A",X"EB23",X"EC05",X"ECF7",X"EDD5",X"EE90",X"EF28",X"EF9C",X"F013",
		X"F0B0",X"F14A",X"F1F2",X"F2C5",X"F3AF",X"F4C2",X"F5EC",X"F6FD",X"F830",X"F921",X"F9EA",X"FAB1",X"FB45",X"FBA6",X"FBEE",X"FC44",
		X"FCAF",X"FD4D",X"FE15",X"FEDC",X"FFB2",X"00B8",X"01C3",X"02BA",X"03E0",X"04D7",X"05D7",X"06AD",X"077C",X"087F",X"0962",X"0A31",
		X"0B07",X"0BB2",X"0C40",X"0CDE",X"0D6D",X"0DFF",X"0E5B",X"0EAE",X"0EDC",X"0EF9",X"0F00",X"0EFE",X"0ED0",X"0E87",X"0E22",X"0DB3",
		X"0D22",X"0CB7",X"0C54",X"0C04",X"0BEB",X"0BE2",X"0C2A",X"0C7F",X"0CFF",X"0D7E",X"0E1D",X"0ECC",X"0F14",X"0F34",X"0F28",X"0F03",
		X"0ED9",X"0EA7",X"0E60",X"0E0D",X"0DB5",X"0D71",X"0D51",X"0D3C",X"0D35",X"0D27",X"0D4E",X"0D62",X"0D6D",X"0D31",X"0CC6",X"0C44",
		X"0BB0",X"0AF1",X"0A16",X"0946",X"0864",X"076A",X"0677",X"059B",X"04B2",X"03E9",X"0327",X"0258",X"019E",X"00C5",X"FFF9",X"FF2B",
		X"FE35",X"FD29",X"FC37",X"FB3E",X"FA41",X"F949",X"F847",X"F736",X"F606",X"F4E6",X"F39B",X"F26C",X"F137",X"EFFB",X"EED5",X"EDD8",
		X"ED28",X"ECBC",X"EC98",X"EC78",X"EC53",X"EC73",X"EC90",X"ECDE",X"ED48",X"ED7C",X"ED97",X"ED9D",X"EDB8",X"EDF4",X"EE1E",X"EE5C",
		X"EE7B",X"EEA3",X"EEEA",X"EF4B",X"EFFC",X"F0A2",X"F16C",X"F248",X"F321",X"F3EE",X"F4B4",X"F584",X"F673",X"F74C",X"F80A",X"F8B9",
		X"F975",X"FA65",X"FB53",X"FC62",X"FD76",X"FE5B",X"FF21",X"FFD0",X"0048",X"00B1",X"00D6",X"00C1",X"00C9",X"00AD",X"00B7",X"00F4",
		X"013D",X"01B7",X"0240",X"02F2",X"03FC",X"0519",X"061C",X"0727",X"07E5",X"0881",X"092B",X"09B8",X"0A3D",X"0AD1",X"0B7F",X"0C21",
		X"0CD2",X"0DBB",X"0E9B",X"0F55",X"0FF7",X"1054",X"1084",X"1077",X"1035",X"100B",X"0FCB",X"0F64",X"0EFB",X"0E80",X"0E0E",X"0DAB",
		X"0D6B",X"0D51",X"0D3D",X"0D18",X"0D00",X"0CEC",X"0CF3",X"0CFF",X"0D16",X"0D16",X"0CFE",X"0CDF",X"0C95",X"0C7C",X"0C57",X"0C03",
		X"0B8A",X"0AEE",X"0A11",X"093D",X"0853",X"0757",X"063C",X"04FE",X"03E6",X"02A5",X"0147",X"0024",X"FF07",X"FDF5",X"FD0F",X"FBEF",
		X"FAFA",X"FA0F",X"F902",X"F832",X"F757",X"F69C",X"F5F8",X"F567",X"F52C",X"F521",X"F510",X"F539",X"F538",X"F510",X"F4C7",X"F442",
		X"F3E1",X"F335",X"F267",X"F18C",X"F094",X"EFBB",X"EF33",X"EEB7",X"EE69",X"EE52",X"EE43",X"EE82",X"EF0A",X"EFA2",X"F04B",X"F0E4",
		X"F186",X"F226",X"F2C7",X"F398",X"F466",X"F50F",X"F5AD",X"F658",X"F722",X"F825",X"F944",X"FA2C",X"FAD6",X"FB67",X"FBA4",X"FB9F",
		X"FBA9",X"FB70",X"FB21",X"FABD",X"FA64",X"FA69",X"FA94",X"FAFF",X"FBD0",X"FCDF",X"FDF4",X"FF41",X"0087",X"01BF",X"02E5",X"03E0",
		X"04AD",X"054E",X"05D4",X"064D",X"06AB",X"0719",X"07B7",X"0835",X"089E",X"0931",X"09AA",X"0A0B",X"0A2A",X"0A39",X"0A10",X"0982",
		X"091B",X"0874",X"07E4",X"0771",X"06D8",X"0691",X"0645",X"060A",X"062F",X"0643",X"0648",X"0661",X"067B",X"06C6",X"0717",X"0765",
		X"07B9",X"0821",X"08A0",X"0916",X"098D",X"0A07",X"0A7B",X"0AE5",X"0B29",X"0B2C",X"0B02",X"0A89",X"09FB",X"0970",X"08DB",X"0845",
		X"0784",X"06B5",X"0610",X"0573",X"04FB",X"049F",X"045F",X"0404",X"03CE",X"0399",X"0392",X"0374",X"035A",X"0341",X"0319",X"02F8",
		X"0290",X"024C",X"0204",X"019F",X"013A",X"00B7",X"001D",X"FFA5",X"FF12",X"FE7C",X"FDEB",X"FD40",X"FC8A",X"FBA2",X"FAC2",X"FA21",
		X"F980",X"F8E4",X"F884",X"F81A",X"F7B0",X"F760",X"F708",X"F6BC",X"F66A",X"F613",X"F5A3",X"F55B",X"F535",X"F4F0",X"F4D1",X"F4DD",
		X"F4E6",X"F515",X"F54D",X"F5A7",X"F5FC",X"F668",X"F6D2",X"F723",X"F78D",X"F808",X"F87E",X"F905",X"F98E",X"FA01",X"FA9D",X"FB33",
		X"FBAA",X"FC1C",X"FC8C",X"FCE6",X"FD34",X"FD99",X"FE0B",X"FE71",X"FEE0",X"FF42",X"FFA7",X"0030",X"00DB",X"0161",X"01F8",X"0264",
		X"02B8",X"02EC",X"02D8",X"02D0",X"0281",X"0239",X"0210",X"01D1",X"01BD",X"01B7",X"0197",X"0191",X"017E",X"0194",X"01C8",X"01BF",
		X"01AA",X"01B6",X"01A8",X"01B9",X"01DF",X"021D",X"025F",X"02B4",X"030E",X"0371",X"03DC",X"042F",X"0487",X"04CC",X"0509",X"0521",
		X"0544",X"053A",X"0531",X"0536",X"051B",X"050D",X"04FE",X"04E3",X"04DD",X"04EA",X"04E9",X"04EA",X"04D0",X"04AF",X"049C",X"0489",
		X"0474",X"047E",X"0488",X"0470",X"048F",X"04B0",X"04D3",X"04D6",X"04D0",X"04D7",X"04F5",X"04FC",X"04FF",X"0501",X"04EC",X"04EB",
		X"04B1",X"0478",X"0440",X"03C0",X"0336",X"0294",X"01D9",X"0135",X"008F",X"FFF2",X"FF6F",X"FEF5",X"FE8F",X"FE3F",X"FDD7",X"FD7F",
		X"FD32",X"FCF0",X"FCE7",X"FCBA",X"FC7B",X"FC58",X"FC24",X"FBE7",X"FBBC",X"FB8C",X"FBA4",X"FB8E",X"FB93",X"FBE9",X"FC18",X"FC48",
		X"FC84",X"FC82",X"FC9C",X"FC68",X"FC29",X"FBE2",X"FB4E",X"FAF8",X"FABB",X"FA42",X"F9A7",X"F941",X"F8E8",X"F8AB",X"F88F",X"F88C",
		X"F888",X"F8AF",X"F8EB",X"F946",X"F9C0",X"FA2B",X"FA89",X"FAC1",X"FAA8",X"FACA",X"FACA",X"FAB2",X"FA9B",X"FA96",X"FAA5",X"FAC0",
		X"FAF6",X"FB69",X"FBA4",X"FBD0",X"FC08",X"FC02",X"FC21",X"FC30",X"FC73",X"FC98",X"FCA1",X"FC95",X"FC9E",X"FC9E",X"FCA9",X"FCC3",
		X"FCE2",X"FD27",X"FD55",X"FDC8",X"FE5B",X"FF00",X"FF9B",X"000C",X"0059",X"00B5",X"0119",X"015C",X"01B1",X"01F2",X"0258",X"02E1",
		X"0385",X"044A",X"0502",X"05C4",X"0688",X"0756",X"0810",X"08C4",X"095C",X"0A04",X"0A9D",X"0AF7",X"0B55",X"0BA5",X"0BF1",X"0C03",
		X"0C13",X"0C01",X"0BC9",X"0B9A",X"0B93",X"0BA8",X"0BC9",X"0BFC",X"0BFA",X"0BD3",X"0BCD",X"0BD1",X"0B8B",X"0B2A",X"0A9D",X"09F7",
		X"094F",X"089D",X"080E",X"0764",X"068D",X"05C8",X"052B",X"048A",X"042A",X"03F5",X"03C7",X"038B",X"0369",X"0374",X"0351",X"030C",
		X"0297",X"0216",X"0175",X"00B4",X"0015",X"FF54",X"FE92",X"FDE4",X"FD2A",X"FC7F",X"FBCE",X"FB13",X"FA54",X"F971",X"F8AB",X"F7D3",
		X"F6C4",X"F5DD",X"F500",X"F427",X"F382",X"F2E8",X"F26C",X"F245",X"F257",X"F2B3",X"F32F",X"F3A3",X"F408",X"F4A0",X"F504",X"F563",
		X"F583",X"F58D",X"F5A1",X"F582",X"F582",X"F56A",X"F565",X"F546",X"F515",X"F50A",X"F522",X"F541",X"F58A",X"F5B3",X"F615",X"F694",
		X"F71F",X"F7DD",X"F87E",X"F923",X"F9E3",X"FA90",X"FB37",X"FBD0",X"FC69",X"FD1B",X"FDAE",X"FE63",X"FEFA",X"FF93",X"0040",X"00BA",
		X"0182",X"0235",X"02B6",X"0347",X"0378",X"03A3",X"0406",X"0457",X"04D2",X"0537",X"056A",X"05CE",X"0600",X"0671",X"06C4",X"06E6",
		X"070A",X"0718",X"073C",X"075E",X"078D",X"07CE",X"0825",X"087D",X"08ED",X"0954",X"09C7",X"0A26",X"0A8A",X"0AFB",X"0B35",X"0B6E",
		X"0B83",X"0B6B",X"0B5E",X"0B22",X"0A99",X"0A3D",X"09BF",X"090C",X"0881",X"07F5",X"0794",X"0746",X"06ED",X"06AD",X"066C",X"062A",
		X"05FC",X"05AA",X"0546",X"04FE",X"0460",X"03E0",X"036E",X"0302",X"02D5",X"02B6",X"028F",X"0274",X"026D",X"0275",X"02B0",X"02AF",
		X"0284",X"0226",X"01C9",X"0157",X"00CC",X"004B",X"FFC7",X"FF55",X"FEEC",X"FEA5",X"FE80",X"FE7A",X"FE83",X"FE88",X"FE98",X"FE79",
		X"FE65",X"FE3F",X"FDD9",X"FD70",X"FD05",X"FC8A",X"FC1E",X"FB98",X"FAF5",X"FA8A",X"FA3E",X"F9C6",X"F966",X"F8E5",X"F86F",X"F7F0",
		X"F785",X"F712",X"F682",X"F612",X"F581",X"F51D",X"F4A5",X"F430",X"F3D2",X"F38D",X"F36B",X"F38F",X"F3A8",X"F3CE",X"F42E",X"F48E",
		X"F4EA",X"F52E",X"F572",X"F5A9",X"F5FA",X"F669",X"F6E9",X"F764",X"F7CC",X"F841",X"F8BF",X"F93D",X"F9B1",X"F9E6",X"F9E6",X"F9EF",
		X"F9CD",X"F9EE",X"FA0C",X"FA3F",X"FAA9",X"FB04",X"FBC0",X"FCBE",X"FDBA",X"FEE4",X"000E",X"0132",X"0228",X"02FC",X"03BA",X"0479",
		X"0508",X"0585",X"05CC",X"0606",X"0684",X"0706",X"07BC",X"0862",X"08EF",X"0966",X"09B1",X"0A0D",X"0A49",X"0A52",X"0A4C",X"0A2F",
		X"0A1D",X"09F7",X"0A22",X"0A61",X"0A9F",X"0AE1",X"0B40",X"0B8F",X"0BD4",X"0BF8",X"0C0C",X"0C21",X"0BF9",X"0BBD",X"0B7A",X"0B3D",
		X"0AE6",X"0A68",X"09FB",X"0961",X"08D6",X"082D",X"0764",X"06D6",X"0606",X"054D",X"04BD",X"03E5",X"031F",X"024F",X"01A0",X"0143",
		X"00D8",X"00A5",X"0085",X"006D",X"0070",X"0068",X"0050",X"0033",X"FFDF",X"FF6B",X"FF00",X"FE76",X"FE05",X"FD9C",X"FD0E",X"FCA3",
		X"FC64",X"FC20",X"FBEE",X"FBB7",X"FB43",X"FADF",X"FA43",X"F9B4",X"F929",X"F892",X"F827",X"F7B0",X"F73C",X"F702",X"F6AF",X"F6A7",
		X"F6AE",X"F69B",X"F6C9",X"F6FF",X"F754",X"F78A",X"F7C9",X"F803",X"F81E",X"F827",X"F81B",X"F7FA",X"F7F2",X"F7B2",X"F782",X"F79A",
		X"F797",X"F798",X"F793",X"F78A",X"F78C",X"F7B3",X"F7B2",X"F7A8",X"F7B5",X"F803",X"F84D",X"F86E",X"F8A0",X"F8E7",X"F947",X"F9D0",
		X"FA70",X"FB1F",X"FBCF",X"FC79",X"FD57",X"FE3E",X"FF22",X"FFF5",X"0099",X"011E",X"01B1",X"022F",X"02AD",X"032E",X"0392",X"03E9",
		X"045C",X"04C0",X"052A",X"058B",X"05E5",X"063F",X"067B",X"06D4",X"0727",X"077A",X"07E2",X"0843",X"0874",X"0893",X"08BA",X"08EC",
		X"0936",X"0944",X"0952",X"097D",X"0999",X"09CB",X"0A02",X"0A48",X"0AA2",X"0ACD",X"0AE9",X"0AF0",X"0AD8",X"0AAF",X"0A52",X"09E2",
		X"0985",X"090E",X"08A1",X"084E",X"0817",X"07F1",X"07D7",X"07D4",X"07B1",X"0792",X"077B",X"076A",X"072A",X"06CA",X"065A",X"05D9",
		X"0573",X"04EC",X"044F",X"03A1",X"02CE",X"0230",X"01BA",X"0150",X"00CB",X"003F",X"FFB4",X"FF3F",X"FEC5",X"FE5F",X"FDEE",X"FD6D",
		X"FCFD",X"FC6E",X"FC2A",X"FBE6",X"FB75",X"FB1C",X"FAD0",X"FA80",X"FA40",X"F9F5",X"F9B2",X"F98A",X"F925",X"F8CD",X"F87D",X"F809",
		X"F77C",X"F6D6",X"F659",X"F5D4",X"F56C",X"F52A",X"F4F6",X"F4CE",X"F4C3",X"F4CB",X"F4EC",X"F528",X"F55F",X"F5A4",X"F5CF",X"F60D",
		X"F652",X"F68D",X"F6C9",X"F707",X"F75E",X"F787",X"F7C6",X"F83D",X"F8BB",X"F927",X"F9A8",X"FA44",X"FAD3",X"FB43",X"FBCE",X"FC6C",
		X"FCDF",X"FD43",X"FDA5",X"FE1A",X"FE66",X"FEC7",X"FF3C",X"FF99",X"0009",X"0075",X"00E1",X"0149",X"01BA",X"0219",X"027A",X"02C0",
		X"02EC",X"0326",X"0351",X"037A",X"0398",X"037D",X"0392",X"03B5",X"03C2",X"03EE",X"0406",X"0427",X"044D",X"0476",X"04B3",X"04F6",
		X"0543",X"0590",X"05C4",X"05FF",X"061D",X"0629",X"061A",X"062C",X"0621",X"05F7",X"05E3",X"05D3",X"05E2",X"05F7",X"0601",X"0610",
		X"062E",X"0643",X"0655",X"0650",X"0643",X"0635",X"0602",X"05C9",X"05AB",X"059E",X"056A",X"052F",X"050C",X"04E9",X"04E6",X"04D3",
		X"04D4",X"04C3",X"04AC",X"04CC",X"04E1",X"04D8",X"04C7",X"048E",X"0476",X"044D",X"0430",X"03EE",X"0394",X"031F",X"02B1",X"0257",
		X"01FE",X"01C1",X"0175",X"0123",X"010B",X"00DD",X"0083",X"002C",X"FFB2",X"FF4A",X"FEC6",X"FE52",X"FDBF",X"FD24",X"FCA6",X"FC58",
		X"FC01",X"FBB2",X"FB66",X"FB19",X"FADB",X"FAA9",X"FA5D",X"FA32",X"F9CB",X"F968",X"F91E",X"F8E4",X"F8B0",X"F85F",X"F83C",X"F821",
		X"F7FF",X"F7DA",X"F7E2",X"F7B5",X"F776",X"F73F",X"F710",X"F70D",X"F715",X"F700",X"F708",X"F728",X"F740",X"F76F",X"F791",X"F79E",
		X"F78E",X"F78F",X"F79A",X"F785",X"F7A7",X"F7B6",X"F7D9",X"F80A",X"F82B",X"F87B",X"F8E8",X"F94C",X"F989",X"F9E1",X"FA3D",X"FAAE",
		X"FB23",X"FBA1",X"FC26",X"FC95",X"FD2A",X"FD9F",X"FE2A",X"FECB",X"FF78",X"FFF4",X"0083",X"0137",X"01C1",X"025E",X"02E1",X"038F",
		X"040A",X"047C",X"04D7",X"054F",X"05CE",X"062E",X"06A3",X"0706",X"0766",X"0799",X"07FF",X"085A",X"08A6",X"08E1",X"0912",X"0943",
		X"0989",X"09CF",X"0A1E",X"0A59",X"0A89",X"0ACA",X"0AFD",X"0B21",X"0B52",X"0B55",X"0B2D",X"0B1A",X"0B14",X"0B1E",X"0B28",X"0B27",
		X"0B31",X"0B24",X"0AF5",X"0ACF",X"0A9B",X"0A5E",X"0A09",X"09A9",X"0954",X"0919",X"08C6",X"089C",X"0882",X"0854",X"0802",X"07A8",
		X"0754",X"06E4",X"0667",X"05BF",X"04F1",X"0431",X"0382",X"02B9",X"01F6",X"0140",X"0073",X"FFD5",X"FF0F",X"FE48",X"FDBE",X"FD1F",
		X"FC94",X"FC15",X"FBA1",X"FB2D",X"FAB7",X"FA4F",X"FA0A",X"F9D0",X"F962",X"F8FE",X"F86A",X"F7FF",X"F7B7",X"F743",X"F6E0",X"F683",
		X"F644",X"F607",X"F5D8",X"F5B5",X"F582",X"F558",X"F53D",X"F53A",X"F52C",X"F52D",X"F50B",X"F509",X"F4E8",X"F4D4",X"F4DD",X"F4CB",
		X"F4D7",X"F4D4",X"F4F0",X"F519",X"F546",X"F568",X"F565",X"F566",X"F58C",X"F5AF",X"F5C2",X"F5BF",X"F5A1",X"F5AC",X"F611",X"F690",
		X"F6FF",X"F76C",X"F7F7",X"F870",X"F922",X"F9C7",X"FA53",X"FAD7",X"FB47",X"FBD4",X"FC50",X"FCB3",X"FD1E",X"FD84",X"FDF3",X"FE7A",
		X"FF01",X"FF92",X"002E",X"00B0",X"0158",X"0214",X"02AF",X"0348",X"03D7",X"0472",X"0545",X"0613",X"069B",X"070D",X"0783",X"07FC",
		X"088D",X"092C",X"09AD",X"0A21",X"0A51",X"0A97",X"0AE8",X"0B23",X"0B7B",X"0BBA",X"0BEC",X"0C26",X"0C70",X"0CB9",X"0CF8",X"0D26",
		X"0D27",X"0D1D",X"0D0C",X"0CF3",X"0CE5",X"0CBC",X"0C95",X"0C73",X"0C40",X"0C2B",X"0C17",X"0C05",X"0BFC",X"0BB9",X"0B6A",X"0B07",
		X"0A7C",X"09F7",X"095E",X"08B5",X"0830",X"0791",X"0703",X"0698",X"062D",X"05D9",X"059F",X"0538",X"04AF",X"043D",X"03A9",X"032C",
		X"0264",X"0194",X"00D4",X"FFE6",X"FF0E",X"FE4F",X"FD9F",X"FCEE",X"FC5A",X"FBDA",X"FB4E",X"FADB",X"FA77",X"FA18",X"F9AA",X"F928",
		X"F86F",X"F7ED",X"F750",X"F6DC",X"F653",X"F5C1",X"F547",X"F502",X"F4A5",X"F45C",X"F430",X"F3F7",X"F3E9",X"F3CC",X"F3B0",X"F374",
		X"F379",X"F35C",X"F358",X"F366",X"F370",X"F360",X"F37E",X"F375",X"F388",X"F3A6",X"F3D2",X"F40F",X"F446",X"F4AE",X"F504",X"F575",
		X"F5CF",X"F634",X"F69B",X"F6E9",X"F734",X"F78C",X"F801",X"F856",X"F8C5",X"F930",X"F998",X"FA28",X"FAC1",X"FB6D",X"FBE3",X"FC61",
		X"FCE6",X"FD85",X"FE21",X"FED1",X"FF6B",X"FFF7",X"007C",X"00F4",X"016B",X"01E1",X"024A",X"02C3",X"036F",X"03EC",X"048E",X"0515",
		X"05AD",X"065A",X"06CA",X"073B",X"07AC",X"07E5",X"0849",X"08AA",X"0910",X"097C",X"09D1",X"0A35",X"0A9B",X"0B08",X"0B7F",X"0BD9",
		X"0BE0",X"0BF0",X"0C1D",X"0C32",X"0C23",X"0C1F",X"0C19",X"0BF7",X"0BEB",X"0BE6",X"0BDF",X"0BD1",X"0B89",X"0B57",X"0B20",X"0AEC",
		X"0AA0",X"0A4D",X"09F2",X"097D",X"08FC",X"0892",X"0819",X"07B2",X"0748",X"06C0",X"066D",X"05E6",X"056E",X"04FA",X"048A",X"040A",
		X"0385",X"0324",X"02CC",X"0261",X"01F3",X"0187",X"011B",X"00D2",X"0050",X"FFE3",X"FF9D",X"FF2F",X"FEB6",X"FE24",X"FD9B",X"FD3C",
		X"FCC9",X"FC57",X"FBC3",X"FB5C",X"FADC",X"FA58",X"F9E6",X"F962",X"F8F3",X"F886",X"F826",X"F7D3",X"F79A",X"F761",X"F735",X"F6FD",
		X"F6CD",X"F68A",X"F648",X"F60E",X"F5C9",X"F58E",X"F56F",X"F547",X"F509",X"F4EA",X"F4CF",X"F4C4",X"F4C5",X"F4C4",X"F4CF",X"F50C",
		X"F546",X"F56E",X"F5A1",X"F5E0",X"F632",X"F6A4",X"F70C",X"F74E",X"F79D",X"F7F3",X"F84D",X"F8A2",X"F8EF",X"F94D",X"F9AE",X"FA0A",
		X"FA9E",X"FB33",X"FBDA",X"FC5F",X"FCE0",X"FD7E",X"FE10",X"FE8F",X"FF25",X"FFAF",X"0010",X"008A",X"00F7",X"017B",X"020D",X"0296",
		X"0310",X"037E",X"03E8",X"0459",X"04D3",X"053C",X"05A1",X"05E6",X"0620",X"0677",X"06D4",X"0738",X"0777",X"07B5",X"07EC",X"0843",
		X"08A3",X"08F7",X"093C",X"0975",X"0988",X"0999",X"09D3",X"0A05",X"0A1B",X"0A2B",X"0A1E",X"0A32",X"0A2D",X"0A23",X"0A26",X"0A26",
		X"0A16",X"09F4",X"09CA",X"096D",X"0930",X"08D5",X"0876",X"0800",X"078F",X"0713",X"06C3",X"067B",X"0633",X"05D8",X"0558",X"04F3",
		X"0487",X"041F",X"03D7",X"035D",X"02E8",X"0251",X"01B3",X"0140",X"00D1",X"0070",X"FFF5",X"FF7C",X"FF1B",X"FECD",X"FE6A",X"FE2B",
		X"FDD7",X"FD76",X"FD3D",X"FCF2",X"FC9E",X"FC69",X"FC1F",X"FBC9",X"FB82",X"FB3C",X"FAFF",X"FABE",X"FA7F",X"FA62",X"FA3F",X"FA0C",
		X"F9D3",X"F996",X"F965",X"F932",X"F8EE",X"F8B6",X"F88F",X"F85F",X"F841",X"F826",X"F818",X"F808",X"F804",X"F805",X"F80C",X"F803",
		X"F7EB",X"F7ED",X"F80B",X"F846",X"F853",X"F871",X"F898",X"F8C7",X"F909",X"F952",X"F979",X"F9B1",X"F9CD",X"F9F8",X"FA6D",X"FAC6",
		X"FB01",X"FB55",X"FB99",X"FBD7",X"FC0E",X"FC4A",X"FCA0",X"FCD7",X"FD0C",X"FD4F",X"FD90",X"FDC5",X"FE36",X"FEA8",X"FF11",X"FF8D",
		X"FFF3",X"0038",X"0073",X"00C7",X"0136",X"0189",X"01CC",X"01F4",X"021C",X"0249",X"0292",X"02E4",X"0303",X"0323",X"0326",X"035E",
		X"03A6",X"03EC",X"0435",X"0450",X"0461",X"0487",X"04D9",X"0517",X"053B",X"0542",X"054A",X"057D",X"05A8",X"05D4",X"05FD",X"0619",
		X"0628",X"062A",X"061B",X"060C",X"05E1",X"05C2",X"05B8",X"0580",X"055E",X"055D",X"057C",X"0584",X"0593",X"059C",X"059C",X"05A5",
		X"05A5",X"0589",X"0547",X"050F",X"04AF",X"0460",X"0414",X"03C5",X"0360",X"0309",X"02D1",X"0298",X"0277",X"0263",X"024B",X"021D",
		X"0210",X"01FD",X"01E0",X"01A2",X"0166",X"0120",X"00CC",X"006B",X"FFF2",X"FFA3",X"FF52",X"FF01",X"FEE8",X"FEAB",X"FE69",X"FE3D",
		X"FE12",X"FE1B",X"FE06",X"FDDC",X"FDA7",X"FD90",X"FD94",X"FD8E",X"FD6C",X"FD35",X"FD21",X"FD1B",X"FD1A",X"FCFF",X"FCC3",X"FC7C",
		X"FC6B",X"FC37",X"FC20",X"FC01",X"FBC0",X"FBB7",X"FBA1",X"FB90",X"FB97",X"FB9A",X"FB9C",X"FBB9",X"FBCE",X"FBDD",X"FBE9",X"FBF5",
		X"FC22",X"FC3F",X"FC57",X"FC69",X"FC7D",X"FC77",X"FC73",X"FC5F",X"FC3D",X"FC25",X"FC29",X"FC36",X"FC4B",X"FC99",X"FCC0",X"FCDA",
		X"FD1A",X"FD89",X"FDDD",X"FE4F",X"FE85",X"FEC6",X"FEDB",X"FF06",X"FF51",X"FF65",X"FF6A",X"FF56",X"FF58",X"FF68",X"FF77",X"FF9A",
		X"FFBB",X"FFC9",X"000A",X"0053",X"009F",X"00D1",X"00DD",X"0107",X"0112",X"013B",X"015D",X"015B",X"017D",X"01A4",X"01D7",X"01EE",
		X"0213",X"0240",X"0272",X"02B5",X"0305",X"031A",X"032A",X"034C",X"0361",X"0384",X"03A3",X"0395",X"0380",X"035A",X"0330",X"031B",
		X"0329",X"0348",X"035B",X"0368",X"0385",X"0397",X"03A7",X"03AA",X"0393",X"038D",X"0367",X"0357",X"0342",X"0315",X"02EB",X"02C8",
		X"02CB",X"02DC",X"02D3",X"02CB",X"02A1",X"0281",X"025F",X"0226",X"0202",X"01BA",X"015C",X"012E",X"00E9",X"00B6",X"0055",X"0011",
		X"000F",X"000D",X"0003",X"FFDE",X"FFD2",X"FFBD",X"FFCB",X"FFED",X"FFD8",X"FF8F",X"FF77",X"FF53",X"FF44",X"FF1D",X"FEE8",X"FEB1",
		X"FE84",X"FE48",X"FE38",X"FE15",X"FDEA",X"FDC4",X"FDAA",X"FDA6",X"FDA8",X"FD9B",X"FD84",X"FD75",X"FD67",X"FD62",X"FD48",X"FD3E",
		X"FD0D",X"FCCE",X"FCB8",X"FCB5",X"FCC1",X"FCEA",X"FCE4",X"FCF4",X"FD08",X"FD00",X"FCEF",X"FCE7",X"FCD0",X"FCCD",X"FCCE",X"FCD3",
		X"FCE2",X"FCDC",X"FCD8",X"FCEA",X"FD0C",X"FD35",X"FD62",X"FD6D",X"FD76",X"FD80",X"FD77",X"FD9A",X"FDBC",X"FDD9",X"FDFE",X"FE1F",
		X"FE46",X"FE64",X"FEB0",X"FEE2",X"FF35",X"FF79",X"FFAA",X"FFEF",X"0019",X"005B",X"0085",X"00C7",X"00F8",X"011F",X"014F",X"0177",
		X"01C1",X"01F0",X"020D",X"0232",X"0286",X"02B0",X"02C6",X"02F6",X"0320",X"0318",X"033F",X"034C",X"032D",X"0338",X"0340",X"032C",
		X"0320",X"0317",X"02E9",X"02F0",X"02F1",X"0311",X"030C",X"0315",X"030B",X"0316",X"032A",X"033B",X"0321",X"0315",X"02FD",X"02D2",
		X"02D2",X"02B2",X"0278",X"0239",X"0219",X"01E4",X"019F",X"0169",X"013B",X"00EA",X"00AB",X"0062",X"0019",X"FFFE",X"FFDB",X"FFBD",
		X"FF9F",X"FF9D",X"FFAD",X"FFB6",X"FFA9",X"FFCA",X"FFB9",X"FFB1",X"FFCB",X"FFD7",X"FFA4",X"FF76",X"FF54",X"FF41",X"FF29",X"FF1A",
		X"FEFF",X"FEE8",X"FEEC",X"FEDE",X"FEFC",X"FEEC",X"FED4",X"FEBA",X"FE9C",X"FE9F",X"FE9F",X"FE86",X"FE8C",X"FE7E",X"FE95",X"FE6E",
		X"FE5C",X"FE45",X"FE34",X"FE1B",X"FE22",X"FE27",X"FE16",X"FE05",X"FDFD",X"FE04",X"FE17",X"FE1B",X"FE15",X"FE29",X"FE12",X"FE29",
		X"FE46",X"FE5D",X"FE61",X"FE67",X"FE51",X"FE5E",X"FE86",X"FE9B",X"FEB2",X"FEAD",X"FEBD",X"FECA",X"FEF2",X"FF0E",X"FF1B",X"FF2D",
		X"FF4D",X"FF67",X"FFA9",X"FFDE",X"FFEE",X"0013",X"0028",X"0065",X"0088",X"00B5",X"00B6",X"00C4",X"00DF",X"00FC",X"0104",X"00ED",
		X"00F0",X"0113",X"0136",X"0160",X"014A",X"0132",X"013F",X"016F",X"01AE",X"01D9",X"01E8",X"01F0",X"020E",X"0234",X"0249",X"0257",
		X"0244",X"023A",X"024A",X"025F",X"0279",X"0250",X"0241",X"0256",X"0272",X"0284",X"0286",X"026F",X"0240",X"0231",X"0223",X"01FC",
		X"01BD",X"0180",X"0156",X"011F",X"0112",X"00F6",X"00F3",X"00AC",X"0089",X"0069",X"004B",X"0022",X"FFD8",X"FFA5",X"FF68",X"FF49",
		X"FF3C",X"FF31",X"FEFE",X"FEC4",X"FEA1",X"FE9E",X"FE96",X"FE66",X"FE48",X"FE2B",X"FE19",X"FE0C",X"FE07",X"FE1E",X"FE24",X"FE26",
		X"FE36",X"FE34",X"FE1B",X"FE15",X"FDF0",X"FDF9",X"FE17",X"FE0F",X"FDFE",X"FE1A",X"FE35",X"FE43",X"FE69",X"FE76",X"FE7A",X"FE77",
		X"FE90",X"FEA8",X"FE89",X"FE79",X"FE75",X"FE7A",X"FE7A",X"FE6D",X"FE4E",X"FE5B",X"FE71",X"FEA5",X"FECC",X"FEE8",X"FF0F",X"FF45",
		X"FF64",X"FF6D",X"FF8B",X"FF6B",X"FF5C",X"FF4E",X"FF5E",X"FF63",X"FF65",X"FF90",X"FFB2",X"FFCE",X"FFFA",X"000B",X"002D",X"0043",
		X"0059",X"0087",X"0098",X"0092",X"00A0",X"00BA",X"00BF",X"00C9",X"00CE",X"00D8",X"00D0",X"00E6",X"00ED",X"0105",X"0122",X"0130",
		X"014E",X"0146",X"014A",X"016B",X"0183",X"018F",X"01A6",X"01AE",X"01B0",X"019D",X"019F",X"01AC",X"01C8",X"01C0",X"01BA",X"01C0",
		X"01A6",X"01AB",X"01AB",X"01CE",X"01DA",X"01CC",X"01C3",X"019F",X"01A0",X"01A4",X"019A",X"0174",X"0156",X"0136",X"0129",X"0144",
		X"012D",X"00F0",X"00A4",X"0092",X"007D",X"0060",X"0022",X"0011",X"FFFF",X"FFF8",X"FFFF",X"FFF5",X"FFDC",X"FFCE",X"FFDD",X"FFB0",
		X"FFA5",X"FFA0",X"FFAE",X"FFA7",X"FFBE",X"FFBE",X"FFB2",X"FFB2",X"FF9D",X"FF7D",X"FF5E",X"FF2E",X"FF1A",X"FF04",X"FEF1",X"FEF1",
		X"FEC7",X"FED0",X"FEE7",X"FF16",X"FF56",X"FF75",X"FF8E",X"FFA0",X"FF96",X"FFA7",X"FF97",X"FF96",X"FF6D",X"FF4A",X"FF1E",X"FF00",
		X"FEFA",X"FEE7",X"FED9",X"FE91",X"FE51",X"FE1E",X"FDFC",X"FDFC",X"FE0F",X"FE01",X"FE0E",X"FE20",X"FE4B",X"FE80",X"FEBE",X"FEF6",
		X"FF29",X"FF2B",X"FF2A",X"FF35",X"FF6C",X"FF7D",X"FF69",X"FF67",X"FF6F",X"FF8D",X"FF93",X"FFA2",X"FF9A",X"FF87",X"FF68",X"FF73",
		X"FF7C",X"FFB4",X"FFE8",X"FFF7",X"0004",X"002B",X"005E",X"0096",X"009C",X"00B8",X"00DA",X"00B4",X"00B0",X"0093",X"00A9",X"00CC",
		X"00BE",X"00D6",X"00D3",X"00F1",X"00FE",X"0117",X"0126",X"0126",X"0119",X"00E7",X"00C5",X"00C4",X"00DF",X"00F4",X"00FD",X"00E2",
		X"00F8",X"0107",X"0137",X"013A",X"0125",X"0113",X"010E",X"0134",X"012A",X"010E",X"0103",X"00F3",X"00FA",X"0102",X"011B",X"011B",
		X"00F4",X"00F1",X"00FA",X"00DB",X"00C9",X"00B4",X"009F",X"0098",X"0086",X"0064",X"003C",X"0033",X"0025",X"001A",X"FFF3",X"FFC4",
		X"FF9C",X"FF7E",X"FF67",X"FF77",X"FF9B",X"FFB2",X"FFB7",X"FFD3",X"FFD0",X"FFC0",X"FFAE",X"FFAE",X"FFBF",X"FFA3",X"FF91",X"FF6C",
		X"FF48",X"FF56",X"FF7B",X"FFA1",X"FFA8",X"FFA3",X"FFA6",X"FF8B",X"FF85",X"FF93",X"FF6E",X"FF5A",X"FF36",X"FF09",X"FF29",X"FF37",
		X"FF3F",X"FF33",X"FF07",X"FF0F",X"FF04",X"FF0D",X"FEFE",X"FF03",X"FF22",X"FF46",X"FF4D",X"FF3C",X"FF3D",X"FF5A",X"FF7D",X"FF78",
		X"FF69",X"FF58",X"FF63",X"FF9C",X"FFD1",X"000D",X"0026",X"0028",X"004C",X"006D",X"0059",X"0064",X"006C",X"0050",X"0022",X"0008",
		X"001E",X"000F",X"FFE3",X"FFDF",X"001C",X"0041",X"0073",X"0064",X"007E",X"0099",X"00C0",X"00D9",X"00CE",X"00D1",X"00EF",X"00F3",
		X"00F4",X"00CF",X"00AE",X"00AB",X"00A1",X"008C",X"0087",X"007F",X"006A",X"005B",X"004D",X"0051",X"0050",X"0020",X"FFF7",X"001B",
		X"0034",X"001C",X"0000",X"FFF0",X"FFEA",X"FFF1",X"FFE8",X"FFD6",X"FFC5",X"FFA8",X"FF8F",X"FFB2",X"FFAD",X"FFC3",X"FFBC",X"FFD4",
		X"FFCF",X"FFCC",X"FFD8",X"FFEF",X"0002",X"0001",X"FFEE",X"FFEB",X"0008",X"000C",X"0021",X"0011",X"000C",X"000C",X"0003",X"FFFC",
		X"FFEC",X"FFFC",X"FFF6",X"FFE7",X"FFEE",X"FFF5",X"0016",X"0037",X"0046",X"0039",X"0036",X"0052",X"005C",X"0041",X"0017",X"0009",
		X"FFE4",X"FFCD",X"FFC5",X"FFA4",X"FF9C",X"FF9C",X"FFAA",X"FFA5",X"FF99",X"FF85",X"FF7E",X"FF51",X"FF48",X"FF37",X"FF1A",X"FF22",
		X"FF13",X"FF1D",X"FF3D",X"FF65",X"FF6E",X"FF6F",X"FF9B",X"FFDB",X"FFE3",X"FFE0",X"FFBE",X"FFD1",X"FFE6",X"FFC0",X"FF95",X"FF4F",
		X"FF4B",X"FF6D",X"FF61",X"FF4F",X"FF4D",X"FF5F",X"FF80",X"FFA8",X"FFB7",X"FFE0",X"FFCE",X"FFF0",X"0014",X"0045",X"0060",X"0074",
		X"0051",X"0395",X"05AE",X"049E",X"04A2",X"0436",X"049B",X"0408",X"0369",X"028F",X"01F9",X"01D1",X"01C4",X"01C5",X"0143",X"00D3",
		X"00C7",X"00A4",X"00AE",X"0082",X"008B",X"0092",X"00F4",X"00EA",X"010D",X"004C",X"FFCA",X"0006",X"004C",X"00FA",X"00EA",X"00B0",
		X"00ED",X"00FA",X"0150",X"013C",X"0130",X"00E6",X"00D7",X"00E0",X"0026",X"FE54",X"FD6C",X"FC38",X"F957",X"F757",X"F4F2",X"F311",
		X"F25A",X"F3A2",X"F5A3",X"F80F",X"FBD6",X"FE0A",X"00BE",X"0604",X"098A",X"0A89",X"0934",X"062D",X"0462",X"04D4",X"0501",X"017C",
		X"FAE0",X"F83E",X"FBDA",X"009A",X"03CB",X"03EA",X"03DD",X"02EE",X"05E8",X"09B6",X"077D",X"04A8",X"01D4",X"0068",X"FC68",X"F79C",
		X"F7D5",X"FB64",X"FBF3",X"FDAA",X"0186",X"02FD",X"0649",X"06EE",X"0C5E",X"07EE",X"0288",X"036F",X"FCB0",X"F767",X"F683",X"F6B9",
		X"F596",X"F699",X"FC28",X"0286",X"0409",X"09D2",X"0B44",X"05AC",X"095E",X"0637",X"0372",X"FB84",X"F204",X"EC9F",X"E551",X"EA7F",
		X"F0BA",X"F2A6",X"F541",X"FB54",X"FC6E",X"027F",X"0834",X"0BE6",X"0704",X"002D",X"03C4",X"00A7",X"F867",X"F7A3",X"F5C3",X"F292",
		X"F317",X"FD16",X"0472",X"FBFC",X"F99D",X"034F",X"068F",X"065D",X"0DD3",X"0DA6",X"FD94",X"F62F",X"06E7",X"0CE5",X"0466",X"031F",
		X"08A6",X"00E0",X"F5EE",X"014F",X"0A98",X"01C8",X"FEE0",X"01F7",X"020D",X"F6FF",X"FD8A",X"15AE",X"11F6",X"0C64",X"107E",X"1221",
		X"09DF",X"09E2",X"0DA9",X"0BDB",X"F6D2",X"EF9C",X"FC35",X"FD29",X"019B",X"075C",X"10D0",X"1006",X"13BA",X"23A3",X"275E",X"1594",
		X"0700",X"0148",X"FB23",X"F277",X"EF5F",X"ED9B",X"E58E",X"DDFF",X"EBF4",X"FECA",X"0801",X"15E9",X"14F3",X"0F06",X"011C",X"0904",
		X"0F77",X"00F0",X"F496",X"EA35",X"E809",X"E365",X"EA0D",X"F7B3",X"FEBE",X"FA97",X"04CE",X"0337",X"FC7E",X"FD78",X"03B8",X"030A",
		X"EFFB",X"ECE1",X"EB10",X"E037",X"E771",X"FCEC",X"0666",X"02F9",X"0C1B",X"150A",X"13AA",X"11A7",X"195F",X"10C9",X"FB48",X"F858",
		X"F390",X"EA79",X"E4B3",X"ECC7",X"F8B0",X"F909",X"0430",X"0DD5",X"0993",X"0ED9",X"15B1",X"1A83",X"0F7E",X"08E8",X"0EBC",X"FE75",
		X"F01A",X"F835",X"F92B",X"F7B2",X"F8CC",X"FF89",X"FA84",X"E4DF",X"E8DD",X"F351",X"EA28",X"E5F2",X"E8DE",X"E516",X"D663",X"DA2B",
		X"F334",X"F537",X"F4CF",X"052A",X"0414",X"F8FC",X"FBD6",X"0927",X"0B86",X"FF1C",X"F821",X"EF75",X"E4D7",X"ECA2",X"FFA1",X"0116",
		X"F4C3",X"F70F",X"0C3E",X"0F86",X"0E4F",X"1D30",X"1E3A",X"184A",X"1BE1",X"20B9",X"1248",X"00CB",X"08C2",X"0F93",X"0466",X"0407",
		X"13DD",X"18C1",X"0BD9",X"12C0",X"2AB9",X"24BD",X"1435",X"223E",X"2141",X"0BDC",X"0139",X"1810",X"20AC",X"0977",X"1889",X"207A",
		X"0E67",X"0588",X"1CCF",X"2074",X"03D4",X"FD58",X"0249",X"F14D",X"DD5A",X"EDBE",X"F010",X"DF80",X"E064",X"F80C",X"FAFF",X"E3BC",
		X"F7A0",X"03F1",X"02F1",X"FE91",X"0596",X"FFE4",X"E506",X"EDF2",X"F52E",X"F214",X"E0CD",X"EF5D",X"F210",X"E40C",X"DFA0",X"F7B6",
		X"008E",X"ECFD",X"FCAE",X"F4A6",X"E9D4",X"E21B",X"F104",X"FEE6",X"F0BF",X"FA87",X"05A9",X"FBB0",X"FD12",X"102E",X"1281",X"1682",
		X"107B",X"12AD",X"12DD",X"027B",X"0744",X"FB16",X"FDE3",X"0013",X"F1BC",X"E419",X"E50F",X"F3F2",X"FD0F",X"FBEF",X"025F",X"FD52",
		X"F996",X"064A",X"09FA",X"05FA",X"0850",X"143C",X"17E7",X"0C05",X"0908",X"0BDC",X"02FA",X"07FE",X"0AF5",X"04B5",X"000D",X"F71C",
		X"FDFF",X"085C",X"092E",X"1371",X"06AC",X"02E8",X"083D",X"10F3",X"0CC3",X"055D",X"FE52",X"FDFF",X"FCF3",X"FEE0",X"FD9F",X"F694",
		X"F527",X"F4D9",X"FB41",X"F08A",X"F6B3",X"0156",X"F6A3",X"F32A",X"FD78",X"FDF6",X"F53D",X"EF3A",X"0020",X"F302",X"DC57",X"EAAE",
		X"F579",X"EF2A",X"EF3C",X"F3F5",X"FF1F",X"F6C3",X"F7F0",X"0620",X"FC7E",X"F0B2",X"F144",X"F3AA",X"EEFD",X"EC3C",X"EDE7",X"F0D1",
		X"F13E",X"FFAA",X"0D7A",X"0974",X"F881",X"FF88",X"0759",X"0C6E",X"0C31",X"1A9F",X"2974",X"1859",X"12B7",X"1448",X"282B",X"2A59",
		X"3100",X"315C",X"1DE2",X"1BA9",X"211B",X"1C3E",X"1595",X"11FF",X"17E4",X"13DD",X"0EBD",X"1157",X"0E9A",X"0ED9",X"1CD5",X"1B89",
		X"1317",X"11B3",X"0C4E",X"0754",X"FDE6",X"03A1",X"FC4F",X"F767",X"EE6C",X"F4A2",X"EB6E",X"E29D",X"DBB0",X"DB31",X"E7A1",X"EBB1",
		X"E5F6",X"D219",X"CB47",X"DAAF",X"E868",X"F98E",X"F2B2",X"F31E",X"F6C2",X"FD8E",X"0278",X"0982",X"102B",X"FFC3",X"F4D9",X"F2BB",
		X"F3F2",X"E81E",X"E428",X"DD73",X"DEC2",X"E2CC",X"E4E2",X"EC00",X"EFD8",X"F5EB",X"0446",X"0FB9",X"1DBE",X"1D27",X"22BA",X"2251",
		X"084A",X"081E",X"1630",X"130C",X"0727",X"FFF3",X"FF4B",X"F58D",X"EE82",X"06E2",X"10CA",X"F18C",X"EF92",X"FFDA",X"186C",X"0E6D",
		X"1435",X"1E2A",X"0F44",X"0C96",X"0E6E",X"038C",X"F1A9",X"F5CC",X"FAC6",X"FA25",X"E2F8",X"E4A6",X"E92D",X"EC49",X"EC07",X"E6D3",
		X"E885",X"DFC3",X"E619",X"FC48",X"FC22",X"F890",X"F77D",X"FA6A",X"0607",X"09B0",X"0E3E",X"0D93",X"0540",X"0837",X"0A61",X"FAF2",
		X"F65A",X"EA36",X"EE95",X"F404",X"F81E",X"F234",X"F066",X"0119",X"21C0",X"19D5",X"1EBC",X"2D1A",X"1E76",X"1034",X"1582",X"229D",
		X"1EAB",X"0B5A",X"091A",X"0908",X"FDCA",X"034F",X"0507",X"0851",X"053C",X"0479",X"FB00",X"F7BC",X"0579",X"19B5",X"1FE5",X"1788",
		X"0D96",X"1412",X"080E",X"0B80",X"09DE",X"03EE",X"F347",X"EDCB",X"F0E4",X"FB5B",X"F63A",X"F9D0",X"064C",X"130F",X"1DAC",X"141C",
		X"0C47",X"F8FC",X"FAA3",X"FF29",X"FEBA",X"FF71",X"FC3B",X"EFF1",X"E455",X"EFAE",X"FF59",X"0DF6",X"120F",X"08A9",X"FE06",X"F6B3",
		X"09AC",X"17CE",X"2283",X"1D6A",X"09AF",X"00FD",X"FFF1",X"04D1",X"02D7",X"F861",X"F4DF",X"F77E",X"EBF4",X"EB78",X"EB11",X"E7CA",
		X"E7DA",X"EB26",X"F45F",X"E8DA",X"DADB",X"DAAB",X"D3B4",X"DA8F",X"E916",X"F0BF",X"FCD9",X"F46A",X"EDF7",X"EA00",X"EBFA",X"F2C5",
		X"06C5",X"0D47",X"F74E",X"E4F5",X"ED52",X"F853",X"EFBC",X"F915",X"01C8",X"F70F",X"E76B",X"EBBB",X"00E4",X"F64B",X"0122",X"14C4",
		X"2371",X"12A1",X"0D2E",X"09EF",X"FB48",X"FE38",X"0000",X"F954",X"D607",X"D870",X"DB59",X"DC0E",X"EB6F",X"00F0",X"1372",X"0D67",
		X"0834",X"18B4",X"2CA1",X"331D",X"3217",X"3321",X"25AA",X"1052",X"0B57",X"114B",X"0BD5",X"0BAC",X"0857",X"0262",X"F27F",X"FA00",
		X"FD9B",X"E558",X"E748",X"F8A4",X"09E6",X"0698",X"0A48",X"0D44",X"0563",X"0E21",X"2D92",X"2EBD",X"1CC9",X"13D3",X"0F96",X"0BF3",
		X"0596",X"06D2",X"FDC4",X"F625",X"F37D",X"F7EF",X"FDA1",X"0456",X"0210",X"0827",X"151A",X"1320",X"0937",X"05C2",X"01C7",X"080D",
		X"03C2",X"0153",X"FFAE",X"F968",X"FF5F",X"06DB",X"0D06",X"03C4",X"062A",X"0616",X"028B",X"03F8",X"038C",X"F9FF",X"E605",X"E765",
		X"EB49",X"F7EF",X"EF59",X"F446",X"05A2",X"0E74",X"1409",X"2871",X"2FDE",X"16DD",X"0ED7",X"07EE",X"F628",X"E3B9",X"E758",X"DDE5",
		X"D3F6",X"CFB7",X"ED5D",X"F299",X"EDFA",X"0072",X"17E0",X"1461",X"1208",X"1B23",X"178F",X"F287",X"F867",X"0A99",X"F732",X"DDCE",
		X"D3CA",X"DA4C",X"D3C1",X"E677",X"0189",X"14B7",X"FEED",X"F5CC",X"FE6E",X"06F1",X"FC2C",X"F8A6",X"F24C",X"D1B7",X"B8D3",X"CFF0",
		X"DC87",X"E219",X"E462",X"ECD7",X"F774",X"F687",X"0D57",X"1FC5",X"0E9A",X"FADD",X"F9C9",X"EA45",X"DA42",X"CA8D",X"D83A",X"D5EE",
		X"D2C1",X"D613",X"E241",X"F4A8",X"0433",X"14ED",X"1B4F",X"2140",X"106B",X"0C3D",X"0D2A",X"FFC1",X"FFA8",X"FA6A",X"016F",X"F404",
		X"FD61",X"0A6A",X"0ABF",X"14C0",X"1E56",X"2B8E",X"1A34",X"1FEE",X"2E78",X"34F8",X"344A",X"2080",X"1833",X"1759",X"18B1",X"257A",
		X"267B",X"18EA",X"1171",X"0FAD",X"1C4F",X"28DA",X"1ED5",X"2622",X"1329",X"126B",X"0E7E",X"173C",X"17DA",X"03A4",X"052A",X"0376",
		X"0637",X"01F3",X"15B3",X"0B05",X"FEDF",X"FD87",X"04DA",X"015B",X"EDFA",X"F761",X"EFC1",X"FCC7",X"0ABC",X"1CFB",X"1E21",X"0D86",
		X"08B0",X"1526",X"1E0D",X"15E3",X"1AFE",X"0303",X"02CE",X"08A2",X"0BB5",X"04EB",X"F9CD",X"0413",X"01EA",X"0016",X"FF85",X"F92C",
		X"F1AC",X"F188",X"FA71",X"FA71",X"FC71",X"E9B4",X"E63B",X"E712",X"EE46",X"E228",X"D86C",X"D7B4",X"D78B",X"E726",X"D954",X"E354",
		X"E672",X"D5E5",X"D0F3",X"D3C3",X"E5C3",X"D285",X"CFB4",X"D3F0",X"D983",X"D9E5",X"E190",X"ED43",X"E612",X"E3AD",X"E4EA",X"EFFE",
		X"DE4D",X"D794",X"D8AB",X"D71A",X"D30A",X"D7F7",X"DF37",X"E2DC",X"EFDB",X"012F",X"0D4E",X"1779",X"1491",X"1339",X"18BE",X"2861",
		X"251F",X"2584",X"141D",X"029F",X"FD00",X"F997",X"04E1",X"01E3",X"0659",X"112F",X"1507",X"164B",X"2028",X"2BE4",X"3D98",X"30A3",
		X"2935",X"26FF",X"1F0B",X"14E0",X"116E",X"12F6",X"0C96",X"0609",X"053A",X"0DC6",X"0BF8",X"11ED",X"1322",X"1630",X"1C95",X"1839",
		X"1B7C",X"069B",X"F09C",X"E92F",X"F554",X"FF0C",X"F83B",X"01BE",X"FEFD",X"0239",X"FE0C",X"114B",X"1325",X"0AD8",X"0A1E",X"F61E",
		X"F1BE",X"E277",X"E903",X"F093",X"E9D7",X"E87B",X"E7E4",X"E9D7",X"EB4C",X"0814",X"2051",X"2961",X"1E99",X"28CE",X"2581",X"0B97",
		X"217A",X"263C",X"1270",X"ECA4",X"DB30",X"F0D8",X"EB36",X"EBC4",X"0686",X"0646",X"F0EF",X"0A0B",X"1960",X"1950",X"1132",X"178F",
		X"174C",X"F8D9",X"0D47",X"21F5",X"0E14",X"F5FB",X"EDBF",X"F496",X"0110",X"07CF",X"12B7",X"02C5",X"E015",X"E894",X"F227",X"F37F",
		X"FA84",X"FE91",X"EEF3",X"D3E0",X"EA0A",X"FE65",X"025B",X"07B5",X"0413",X"F4BF",X"E64B",X"F50B",X"07D2",X"01E8",X"FA15",X"0143",
		X"F770",X"E26D",X"F58A",X"0996",X"0246",X"F4FF",X"07AF",X"0E1B",X"ED65",X"FC62",X"1168",X"0E9A",X"013C",X"1338",X"1D34",X"FF30",
		X"057F",X"246A",X"21F6",X"0C31",X"14C4",X"10C0",X"F36E",X"E85C",X"F87D",X"EA76",X"D1C0",X"E0A3",X"E296",X"CE35",X"D297",X"E43B",
		X"F427",X"DD59",X"F3A9",X"FE75",X"E9B7",X"EDFA",X"F21B",X"0198",X"F624",X"F7A8",X"F805",X"E788",X"DE60",X"F774",X"F8EF",X"EB4C",
		X"F2A5",X"F4A9",X"FCF0",X"FA5E",X"0B2A",X"09A9",X"F53E",X"0937",X"0E12",X"F647",X"F35A",X"FD9E",X"FF71",X"F2C5",X"F9C0",X"F928",
		X"E438",X"DE84",X"F163",X"EE26",X"F3F5",X"0D64",X"166E",X"0BF1",X"FF15",X"20E1",X"2C68",X"26EF",X"2F82",X"301A",X"1B60",X"042D",
		X"0114",X"19C1",X"1074",X"FDB7",X"F483",X"EDB5",X"F52B",X"FED1",X"1125",X"02C1",X"F4D8",X"FE52",X"1669",X"108D",X"040D",X"FFE7",
		X"FF6B",X"075A",X"0FAD",X"12E3",X"08B2",X"FF00",X"00FA",X"1AB5",X"163D",X"FE8B",X"05BB",X"14DB",X"113C",X"086D",X"0F77",X"158A",
		X"0EC2",X"1FF6",X"26C0",X"1CEB",X"137D",X"1D34",X"224A",X"1BC2",X"1645",X"1E5A",X"0D89",X"F751",X"0197",X"F54A",X"EDC5",X"E20B",
		X"EEEE",X"F651",X"E3A7",X"F2E2",X"FDFD",X"FD8B",X"0896",X"0B1B",X"0253",X"0C27",X"0980",X"187F",X"143C",X"0D68",X"12B4",X"072E",
		X"0106",X"F098",X"F83A",X"FFA4",X"0576",X"ECA2",X"D7B4",X"C966",X"D914",X"E619",X"E090",X"ED0D",X"E5AB",X"F086",X"13E0",X"1F41",
		X"120F",X"1148",X"10FF",X"0773",X"008F",X"08E2",X"03E4",X"F54A",X"E1E5",X"E548",X"DB43",X"E3E6",X"EA50",X"F267",X"F521",X"F6F8",
		X"02A5",X"0918",X"1565",X"1F0A",X"2E85",X"1688",X"0A01",X"FE78",X"F259",X"E7D6",X"EA42",X"E067",X"CAF5",X"C120",X"CF75",X"DDC8",
		X"DD46",X"E5F3",X"EC8F",X"E939",X"EB4B",X"FA31",X"00D4",X"E2E9",X"E668",X"EEFE",X"E64B",X"DF8A",X"D97D",X"E2E6",X"D65F",X"E24A",
		X"E96C",X"F5B2",X"F732",X"FBDD",X"006E",X"0439",X"12D7",X"1B4D",X"2B48",X"1FE8",X"1BE2",X"18F8",X"1D89",X"1C59",X"12FC",X"0AE5",
		X"05FE",X"FDCD",X"FD45",X"097D",X"03FA",X"FA3B",X"FF38",X"1419",X"2AA7",X"28BE",X"3117",X"349C",X"2271",X"20D5",X"2D59",X"263B",
		X"175F",X"1268",X"0301",X"F815",X"F3BF",X"0CDC",X"1D28",X"08B2",X"0569",X"07AC",X"092B",X"0B5E",X"20F2",X"27BA",X"1028",X"0733",
		X"0789",X"05F7",X"036F",X"0E08",X"0817",X"F731",X"F0DB",X"F961",X"F39D",X"FA1C",X"0E21",X"FC71",X"F46D",X"F3C5",X"04AB",X"FCA0",
		X"E48A",X"D943",X"DD89",X"DBF4",X"E8C4",X"0B1E",X"05D8",X"FD5C",X"FDBD",X"12E0",X"1658",X"1A01",X"2BA1",X"1DAC",X"FE7B",X"FC94",
		X"0E03",X"0085",X"EFD8",X"EDF8",X"F3FF",X"E626",X"DF01",X"FBF2",X"06C8",X"0669",X"122E",X"202E",X"1BA6",X"1506",X"275A",X"2ACD",
		X"14EC",X"11CA",X"115E",X"0DB0",X"F7FF",X"EFD1",X"E502",X"E329",X"DA1E",X"E141",X"F2F8",X"EC85",X"EFE8",X"0743",X"175F",X"0AC5",
		X"1A86",X"2729",X"075C",X"E3D0",X"F9C3",X"0203",X"F2A8",X"EB23",X"F189",X"F414",X"E170",X"F2A6",X"0A5D",X"F28A",X"EDCB",X"FDD0",
		X"FD1F",X"E578",X"ECAE",X"0427",X"E710",X"D1C0",X"E31F",X"EBA8",X"D0FD",X"DCE2",X"DF8E",X"D225",X"C92E",X"E358",X"FA24",X"EACD",
		X"E5DF",X"F454",X"F590",X"E268",X"E218",X"E4F2",X"D523",X"C072",X"D1FA",X"D181",X"B6F2",X"C5EE",X"E4CA",X"EEBE",X"EDAF",X"0230",
		X"16B1",X"02A2",X"0B80",X"1FC6",X"13C1",X"0A37",X"1352",X"1F99",X"0D0C",X"08D1",X"1911",X"18BE",X"08A2",X"1562",X"216D",X"165B",
		X"1A43",X"21F5",X"1BBB",X"0F87",X"234A",X"2F0A",X"2396",X"217D",X"204D",X"1F8F",X"3724",X"4AA3",X"4AF4",X"40A1",X"3D42",X"35BC",
		X"2EEA",X"2D19",X"318D",X"1FF8",X"1536",X"162C",X"142C",X"1B56",X"2318",X"34F1",X"299D",X"262E",X"3321",X"2402",X"1102",X"1CE4",
		X"2362",X"0BF8",X"F8E8",X"018E",X"F37C",X"E64F",X"F9BD",X"FC91",X"E4D9",X"E4E3",X"F5EF",X"F7F5",X"E5FC",X"F017",X"FF8E",X"EBC5",
		X"DBD5",X"E28D",X"E328",X"D31C",X"D572",X"E241",X"D9AB",X"CA7D",X"DFFF",X"F111",X"DD7D",X"D8BE",X"F163",X"F34D",X"E28D",X"DEC3",
		X"E9B5",X"CC9A",X"C7A9",X"E38D",X"E590",X"C8BC",X"CD7B",X"E7C7",X"E335",X"DED8",X"FF05",X"0FA4",X"FE1C",X"0731",X"1B56",X"2451",
		X"1B8E",X"1BB9",X"10C0",X"0252",X"F9D6",X"F935",X"F66A",X"EB7E",X"E335",X"E93F",X"F938",X"014C",X"FD19",X"09D6",X"192D",X"1C49",
		X"200B",X"2E01",X"26A0",X"19FD",X"187B",X"17D7",X"04B5",X"FAD9",X"06E4",X"0210",X"FCBA",X"F58D",X"02A5",X"05E5",X"06AF",X"0D9C",
		X"1792",X"0CFF",X"F747",X"F0B2",X"EAC8",X"E19A",X"D691",X"D689",X"DAB9",X"D2B7",X"BF58",X"C922",X"DB83",X"F0A5",X"F0D5",X"F580",
		X"F0EB",X"E167",X"F7E2",X"159B",X"143F",X"FE2C",X"F94E",X"FD6E",X"F1EB",X"F172",X"0990",X"0CEB",X"0126",X"FD65",X"1D82",X"25B0",
		X"21D9",X"3056",X"3ADF",X"1F99",X"0E27",X"1629",X"0DA3",X"EBCB",X"DD31",X"EA72",X"EB10",X"D9E1",X"EAEC",X"0896",X"00A7",X"13A4",
		X"379A",X"4D84",X"2F9A",X"3269",X"49DE",X"310A",X"0C17",X"1FAF",X"246A",X"0F97",X"FBE9",X"0733",X"138B",X"0459",X"1BB7",X"227D",
		X"1CC1",X"1FEE",X"1E01",X"0C0B",X"00A5",X"0272",X"0DA7",X"FE8B",X"EC33",X"DD6C",X"E435",X"EDB1",X"F6CF",X"EC7F",X"E190",X"DB66",
		X"C979",X"D220",X"E4AA",X"FFFD",X"F7FF",X"E441",X"F0E4",X"FA81",X"0065",X"0550",X"0378",X"ECA1",X"DBCB",X"E1DC",X"F079",X"F27A",
		X"E564",X"E2A3",X"E1E8",X"E47D",X"EA88",X"FCED",X"077D",X"039C",X"060A",X"09AF",X"FF75",X"0E67",X"263A",X"17B1",X"0A18",X"016C",
		X"04CB",X"026C",X"FDCD",X"03F1",X"046F",X"F8BA",X"FC64",X"04D4",X"0AF2",X"0BC8",X"101F",X"12B7",X"0650",X"0D21",X"0C8D",X"0209",
		X"FA29",X"F525",X"F35D",X"FFB1",X"FB0C",X"0272",X"F6E8",X"FDC6",X"1005",X"0A31",X"1015",X"111A",X"09CF",X"08B5",X"0304",X"FF81",
		X"FE64",X"F424",X"FC6C",X"F1AE",X"EA46",X"FF36",X"0677",X"0133",X"FCE0",X"034C",X"1FE6",X"18E1",X"0760",X"078D",X"0566",X"F387",
		X"F2D1",X"E936",X"DC04",X"CD84",X"D11D",X"EDE5",X"F0B5",X"FED4",X"1284",X"21FC",X"21A9",X"2B3F",X"3E0B",X"3C5A",X"2DAA",X"18D2",
		X"0EEB",X"0085",X"E8CC",X"E9C0",X"E53B",X"E16D",X"CEF0",X"D695",X"E85B",X"E858",X"F5E4",X"FDFA",X"0B18",X"F26D",X"EBB8",X"0B60",
		X"06D1",X"FEF3",X"F667",X"F3B6",X"F5C2",X"F18A",X"F3B3",X"06E2",X"FB13",X"FF48",X"082A",X"F56D",X"FDA4",X"0D44",X"2CBE",X"1752",
		X"F341",X"EE85",X"06CE",X"0928",X"11B0",X"0B67",X"05EB",X"02BB",X"FF35",X"2153",X"247A",X"19C8",X"1155",X"09FE",X"0824",X"F9D6",
		X"0053",X"090B",X"F227",X"F764",X"F75E",X"EF8C",X"F011",X"F487",X"FDDA",X"FAC6",X"E20E",X"FBA3",X"F7A7",X"F3BC",X"0B0D",X"0052",
		X"FD54",X"DDAC",X"F657",X"05D4",X"FA1C",X"F2D8",X"E8E0",X"EB37",X"F87D",X"034C",X"EEBF",X"E5D9",X"D10D",X"ED13",X"F289",X"E965",
		X"F45D",X"F2A3",X"061D",X"0BD2",X"1939",X"FF77",X"F8E5",X"F5A6",X"FD52",X"F96B",X"F3E2",X"EEDE",X"DACE",X"EEE1",X"F574",X"00BB",
		X"FDE9",X"00F9",X"0759",X"0953",X"1668",X"278E",X"3386",X"31C8",X"1EB2",X"27DD",X"2E0D",X"226D",X"26D6",X"2D85",X"28E0",X"1E0B",
		X"1C66",X"2E75",X"1B1E",X"1519",X"1F33",X"14D0",X"0E12",X"117E",X"1AFD",X"017C",X"F1B8",X"0D96",X"23D3",X"152F",X"0F37",X"105E",
		X"0C1E",X"F8EF",X"0CC3",X"1071",X"085D",X"E74F",X"F15A",X"00C1",X"FA12",X"FCB8",X"FDF3",X"0546",X"FD48",X"FDD1",X"F658",X"EF82",
		X"E402",X"F2CE",X"F680",X"EC2D",X"E3E0",X"E9AE",X"F2EF",X"FC2B",X"FB5F",X"FE0C",X"0042",X"FA51",X"F77A",X"048B",X"0937",X"FEF3",
		X"F27C",X"F715",X"EC20",X"D703",X"DB04",X"DFDB",X"E1CC",X"CF1F",X"CB08",X"E105",X"E13F",X"D545",X"CF32",X"CD51",X"C489",X"C818",
		X"D976",X"EF50",X"D4A8",X"D76F",X"E419",X"E60C",X"F83E",X"0634",X"FDD7",X"E0E9",X"DA5F",X"F37F",X"F53E",X"E5EC",X"F5A0",X"F2F4",
		X"DB6D",X"D28B",X"ED92",X"FC09",X"F745",X"0192",X"0680",X"FFE4",X"06FB",X"1CE8",X"2D78",X"22F2",X"1FF8",X"147E",X"105E",X"0C7E",
		X"1C79",X"15E0",X"0F71",X"1055",X"1D27",X"22B3",X"10D2",X"0ECC",X"1962",X"1723",X"1707",X"166F",X"03A5",X"010E",X"0CA3",X"2127",
		X"210F",X"1A36",X"1B2A",X"1E60",X"1A50",X"1DD8",X"236B",X"10AB",X"0937",X"0D25",X"16BB",X"0AE2",X"0453",X"01EB",X"0779",X"1439",
		X"2051",X"24F0",X"1E8C",X"2515",X"22E5",X"3537",X"38CC",X"4282",X"3B70",X"2E7E",X"1F93",X"119D",X"0C41",X"0973",X"045F",X"0CB3",
		X"0EC0",X"0138",X"FA38",X"0592",X"0E2E",X"0DD5",X"0268",X"12BA",X"089D",X"FBE9",X"188F",X"18D1",X"1FB5",X"0B86",X"1556",X"0B3D",
		X"F147",X"ED0D",X"0869",X"F921",X"E591",X"DCFB",X"D3E3",X"DDCC",X"D7FA",X"E8D0",X"DBAC",X"CB8A",X"D44B",X"D55F",X"DABE",X"D79E",
		X"D60D",X"ED39",X"ED59",X"F3D2",X"FD42",X"01C8",X"EF52",X"F408",X"F3FB",X"0514",X"038B",X"F9BF",X"F98B",X"F87A",X"FE88",X"F63A",
		X"F2B5",X"F085",X"E45E",X"E603",X"E184",X"CE37",X"CA4A",X"C36C",X"CFFF",X"D258",X"D081",X"C747",X"D536",X"D265",X"DE47",X"F1AC",
		X"04FA",X"04CB",X"FE18",X"0F68",X"FB87",X"F2D2",X"F1E8",X"0761",X"02FD",X"E187",X"DB59",X"E37D",X"EC9E",X"ECDA",X"0200",X"FA15",
		X"EDE4",X"F638",X"FDC9",X"FE9E",X"F641",X"0233",X"F741",X"E9CE",X"ECC1",X"E19D",X"D7A5",X"D349",X"DD11",X"E441",X"F1EE",X"EC13",
		X"FC19",X"FFE1",X"F4B5",X"FCEC",X"02D4",X"0FAD",X"FE55",X"FAD0",X"FCA0",X"FF0D",X"0D38",X"2315",X"28EA",X"27DA",X"2B5B",X"3279",
		X"3341",X"2CA2",X"3B2C",X"4042",X"2FA6",X"230B",X"0E31",X"03B5",X"12D6",X"245A",X"2218",X"1FB9",X"25CA",X"2EBB",X"3DEC",X"4C6A",
		X"5268",X"484D",X"4AE2",X"43BE",X"3099",X"3583",X"3466",X"35EF",X"252B",X"1E3D",X"2502",X"36F4",X"429B",X"2CDE",X"1E25",X"10DA",
		X"1630",X"0B2B",X"19FA",X"1820",X"F899",X"E131",X"EC9B",X"13D6",X"17FD",X"2800",X"2764",X"22C3",X"1D60",X"3C77",X"4B40",X"23FC",
		X"0BEC",X"010A",X"FEF6",X"E389",X"E267",X"E623",X"D5F0",X"D43C",X"EDE0",X"FBC3",X"E914",X"F4FF",X"F9D3",X"F3EB",X"EB59",X"EED1",
		X"E603",X"C269",X"B8CD",X"C023",X"C45A",X"BCFA",X"C94A",X"D1E0",X"D072",X"D2C1",X"EB8B",X"FEE6",X"E4AA",X"E17D",X"EC03",X"E74F",
		X"CC6A",X"C9C9",X"D31F",X"B7F5",X"ABFB",X"BE4B",X"D407",X"C957",X"D798",X"E50F",X"DC64",X"D08A",X"EAED",X"F90F",X"E635",X"D616",
		X"CF38",X"C0BB",X"BB32",X"CEEF",X"DE14",X"DA6D",X"CE74",X"D265",X"E24A",X"EE92",X"EE0A",X"F04D",X"F5E8",X"E4A4",X"DEA3",X"EEFD",
		X"EEDA",X"EEDE",X"ED59",X"01E7",X"09C5",X"02FA",X"0378",X"0CBD",X"0036",X"FDC7",X"FFFD",X"F9A1",X"F67C",X"FF10",X"111F",X"1488",
		X"07C1",X"117E",X"0ED6",X"1B03",X"318D",X"2243",X"17AB",X"0698",X"155F",X"24B9",X"37D6",X"2E4C",X"1F47",X"0F81",X"1235",X"280B",
		X"34FF",X"400A",X"3B1B",X"3F2F",X"33CF",X"323A",X"4162",X"4562",X"3E32",X"30DE",X"263B",X"25B7",X"0D97",X"156B",X"322C",X"33B5",
		X"28FC",X"2B20",X"3753",X"38F8",X"2C5C",X"4620",X"4598",X"2C68",X"3E87",X"303A",X"1814",X"03E8",X"1FA8",X"29B7",X"15E3",X"0130",
		X"117B",X"0F7A",X"08FE",X"1B60",X"260F",X"3192",X"15B7",X"0FE6",X"0D47",X"FFE0",X"F8CC",X"0182",X"F7AA",X"E02D",X"D659",X"E34E",
		X"EA2F",X"EDE1",X"020D",X"110F",X"0137",X"FCA1",X"08B2",X"FA77",X"F280",X"F6D6",X"E94E",X"B577",X"B6D9",X"CB63",X"D4B1",X"C424",
		X"C53D",X"CE4B",X"C3F7",X"DBCB",X"E135",X"EFE5",X"E409",X"DE7A",X"D0E4",X"CF35",X"CE74",X"CC41",X"CB80",X"AC1A",X"A733",X"AB26",
		X"CAAC",X"D55C",X"CDF6",X"CF74",X"C482",X"CA7A",X"D368",X"E8E6",X"EBEA",X"DAFA",X"CBA9",X"C82E",X"C6F7",X"CD3B",X"DD34",X"DD3D",
		X"D139",X"C5E5",X"CF77",X"E5EF",X"EC68",X"F3AC",X"FA2B",X"FE4C",X"F7C3",X"F83B",X"0036",X"FB1F",X"FCD3",X"FF0C",X"05B1",X"FE7E",
		X"0743",X"0D4E",X"0905",X"15CA",X"2221",X"29BD",X"1B2C",X"15B4",X"211C",X"309E",X"3DD3",X"3A6D",X"4032",X"3DA9",X"3BD6",X"3E98",
		X"41A4",X"331A",X"2F11",X"2521",X"1138",X"14A7",X"1377",X"1C4A",X"15DD",X"1CCF",X"23B2",X"2790",X"30D8",X"3818",X"3A1F",X"341E",
		X"3E45",X"34CC",X"2894",X"15B1",X"2264",X"20C6",X"1A17",X"148B",X"0B77",X"0993",X"1B4F",X"3370",X"2928",X"25BC",X"2EEE",X"2B94",
		X"2741",X"2F30",X"3040",X"1C50",X"16A7",X"097D",X"0853",X"076F",X"0880",X"125B",X"0013",X"0807",X"17ED",X"3079",X"2F43",X"1A9C",
		X"1736",X"1D39",X"0695",X"0FA0",X"0840",X"E65B",X"CDC9",X"C96D",X"DF44",X"E93F",X"EE4C",X"F7B0",X"E7E6",X"D84C",X"E8A1",X"04D4",
		X"19B4",X"09D6",X"F6B9",X"E097",X"D65F",X"D970",X"E17D",X"CE2F",X"C072",X"BC49",X"B652",X"D05B",X"CCF9",X"DD8C",X"EDFD",X"F81F",
		X"F044",X"F201",X"F673",X"EDFD",X"E7F7",X"EF70",X"D604",X"BB10",X"C4EB",X"BA8A",X"B5D6",X"AF69",X"CCDF",X"CF47",X"D3C7",X"DAE2",
		X"DD30",X"E4C0",X"DD1E",X"E41B",X"ECBA",X"E1EC",X"D623",X"CE5E",X"CD7A",X"CA70",X"D206",X"D38E",X"E4D6",X"D953",X"CCF9",X"DC14",
		X"E11C",X"F07F",X"F3C5",X"057C",X"04CA",X"F7B6",X"F954",X"F787",X"E833",X"F283",X"FBE9",X"ED50",X"E675",X"DBBF",X"E798",X"EE13",
		X"F20A",X"02C4",X"0DB9",X"05CE",X"FC5B",X"06FE",X"1FF8",X"0F6A",X"18B7",X"2FE4",X"2C13",X"23AD",X"2CA7",X"37D2",X"2E93",X"2E55",
		X"4AD1",X"4CAC",X"301D",X"3DCD",X"510F",X"5568",X"4536",X"46C7",X"4590",X"33D8",X"380C",X"45EE",X"3B48",X"28F6",X"339C",X"3E74",
		X"343A",X"2875",X"2832",X"2D19",X"2102",X"2E7C",X"45FB",X"48A2",X"374A",X"30CE",X"39C6",X"37C6",X"3799",X"42CE",X"329C",X"2180",
		X"1471",X"19D7",X"1588",X"0867",X"18D1",X"0C6D",X"E59E",X"DCC6",X"EEB8",X"F96D",X"F7C9",X"FD7B",X"F94B",X"E7B8",X"E5F3",X"F961",
		X"FB94",X"EF60",X"EF5D",X"EBDE",X"DCB8",X"D6CD",X"DC5B",X"E5B4",X"DFBC",X"E127",X"F1B2",X"EFA6",X"EA5B",X"F8B6",X"04DB",X"0091",
		X"002C",X"0155",X"F276",X"DAEB",X"EBA8",X"EFA8",X"E6D0",X"D579",X"D2F6",X"D17B",X"C495",X"C4BC",X"D67C",X"CB28",X"BF3F",X"C76D",
		X"CE03",X"C19E",X"B0C6",X"BCF6",X"B6E5",X"AD34",X"B044",X"C918",X"C159",X"BBF9",X"CBD5",X"D55F",X"E022",X"E403",X"F635",X"F069",
		X"E4B3",X"E358",X"EC69",X"D9FB",X"CC47",X"D6C1",X"D19D",X"CE6A",X"C715",X"D96F",X"DB0E",X"E75E",X"F02D",X"F428",X"FF29",X"0046",
		X"0F57",X"296B",X"2CC5",X"2AB5",X"2BF0",X"2360",X"23EE",X"1FB3",X"295C",X"2BE3",X"1E96",X"198F",X"177B",X"1497",X"213B",X"31A4",
		X"3560",X"37D9",X"29BA",X"2A52",X"3B18",X"44A5",X"49AF",X"4256",X"40D7",X"2F83",X"2A7C",X"3A51",X"3A7E",X"2F49",X"23DC",X"2645",
		X"25CD",X"14C7",X"1A6F",X"2B55",X"2F1D",X"3AFC",X"2ADA",X"22FB",X"1C2E",X"110A",X"0A44",X"FE8B",X"FA7D",X"FCCA",X"EB66",X"EBB1",
		X"FE84",X"03ED",X"0F86",X"16AD",X"2755",X"2458",X"2597",X"2C89",X"1A8F",X"143F",X"2C4F",X"2247",X"07E8",X"F7F9",X"F211",X"FBB3",
		X"EDAB",X"EAA5",X"F6D6",X"EDF7",X"E9D0",X"FB3B",X"1E61",X"1939",X"1041",X"132C",X"1698",X"0549",X"118E",X"20BF",X"0B89",X"F2CE",
		X"EFCF",X"F752",X"F16C",X"FD28",X"0B6D",X"0B1A",X"F596",X"F844",X"05E7",X"F50B",X"EACE",X"F12D",X"E23B",X"C7EE",X"C7DF",X"D945",
		X"D523",X"CBB3",X"C740",X"C5D7",X"C266",X"D3E4",X"CBF5",X"D1DD",X"D181",X"D194",X"D7CE",X"CADF",X"D005",X"CC87",X"C631",X"C092",
		X"C684",X"C715",X"C07B",X"C4E4",X"D577",X"DF47",X"D403",X"E3A1",X"E51F",X"EBFD",X"E97E",X"EBD7",X"EE03",X"DD5E",X"F5DC",X"F773",
		X"FF72",X"FC67",X"F6B2",X"ED43",X"E209",X"E44F",X"EA6F",X"E0C3",X"D242",X"EC19",X"F460",X"0504",X"0207",X"0776",X"1EF7",X"1B70",
		X"21C2",X"2BBD",X"23CD",X"206D",X"10B0",X"0F3F",X"16E3",X"1781",X"1A24",X"17EA",X"0EA0",X"16EB",X"284F",X"2557",X"2702",X"2B0C",
		X"37FB",X"1D8F",X"12F9",X"14DD",X"0FE5",X"17A1",X"0C4A",X"1044",X"1151",X"0E3F",X"1555",X"19EA",X"3252",X"34A0",X"2BA5",X"3269",
		X"253B",X"1B3A",X"2641",X"293F",X"2056",X"08F5",X"FA84",X"F8B7",X"F9C4",X"103B",X"1DF2",X"1CC1",X"1087",X"17AD",X"2B6F",X"2812",
		X"2CD7",X"3473",X"3958",X"2511",X"233A",X"2F20",X"2512",X"115E",X"0663",X"FB0F",X"F861",X"FAAD",X"FD00",X"F502",X"E874",X"F6B6",
		X"0665",X"070B",X"0E94",X"1E4C",X"1364",X"FC55",X"00C7",X"0336",X"FD46",X"F043",X"ED76",X"F4FB",X"D6E3",X"CD67",X"C5CF",X"C89C",
		X"D8B2",X"E0A9",X"E5A4",X"D5F0",X"CB5A",X"D755",X"E791",X"F176",X"ED9B",X"E212",X"D0E7",X"CA41",X"DD04",X"F36E",X"EF5D",X"E655",
		X"D8A2",X"DAFB",X"D992",X"E985",X"F6CF",X"ED4F",X"EA4C",X"E76B",X"FC05",X"F5BC",X"FA05",X"F3BC",X"E61C",X"E024",X"E38A",X"E5A4",
		X"E5FF",X"E11E",X"ED60",X"E93F",X"EA91",X"020A",X"0BD2",X"1B46",X"035F",X"059F",X"075A",X"05A8",X"1788",X"148F",X"0EE2",X"F42A",
		X"ED8B",X"FFB2",X"FE82",X"F961",X"00A8",X"0BFC",X"04C4",X"F587",X"F7F0",X"FA3B",X"F2A6",X"FDF6",X"F599",X"EFB5",X"E4BA",X"F186",
		X"095C",X"0C5A",X"10E9",X"06BC",X"035F",X"093D",X"1455",X"234E",X"2CFA",X"2747",X"17BE",X"1B2A",X"1A17",X"153C",X"1F7C",X"21A7",
		X"1FDF",X"13AD",X"0EC3",X"140C",X"1409",X"1097",X"109E",X"0EC6",X"097C",X"0B51",X"1C63",X"2FA9",X"2D0A",X"2608",X"2758",X"2FCE",
		X"216C",X"1F8D",X"36F5",X"218E",X"0CCF",X"FF88",X"0CB3",X"0EDC",X"F8D5",X"0CD5",X"0E54",X"0540",X"01C1",X"0E0C",X"2B65",X"2A53",
		X"22BD",X"1ED8",X"1294",X"0989",X"0072",X"0349",X"062D",X"EF00",X"E4C9",X"E0C9",X"DC17",X"E1FC",X"FC0F",X"1A98",X"0250",X"EEDB",
		X"058F",X"2547",X"13D0",X"0DAD",X"14A1",X"F55D",X"DC24",X"D013",X"E358",X"DB8C",X"CA64",X"CC61",X"DAE8",X"DBF8",X"DA1E",X"F461",
		X"F9E9",X"EFD2",X"F8C9",X"0740",X"F9E6",X"E422",X"E134",X"DD1B",X"CC67",X"C77A",X"D6AF",X"CEF0",X"CB8D",X"D701",X"E351",X"D933",
		X"C0C1",X"EB14",X"F90E",X"E32E",X"E22A",X"EB50",X"ED71",X"E54B",X"F286",X"EAEA",X"D507",X"D5E7",X"F1A9",X"EB55",X"E13D",X"E09A",
		X"F9FF",X"F9C0",X"E76B",X"00A7",X"0740",X"F9C5",X"FD5E",X"210D",X"1697",X"F690",X"FF95",X"0449",X"0737",X"11F3",X"22C0",X"23B0",
		X"13F0",X"0BBC",X"196F",X"28E6",X"2DBB",X"2E8B",X"215D",X"18BC",X"19CE",X"208F",X"18FA",X"155C",X"FF00",X"FEBE",X"F8D2",X"03D4",
		X"10AA",X"1CD1",X"3214",X"2597",X"1AFD",X"255B",X"1F5B",X"205E",X"29D3",X"1BD2",X"0743",X"EC76",X"FAD0",X"FC55",X"0191",X"FA32",
		X"F5C2",X"F217",X"FE71",X"0669",X"1BAC",X"1C83",X"15AA",X"0BD6",X"055C",X"00E1",X"0E21",X"202A",X"0F7D",X"FF46",X"FBC0",X"0CFF",
		X"1526",X"250C",X"2651",X"0A5A",X"F2C9",X"FF49",X"0918",X"11FD",X"036C",X"0216",X"EBBB",X"E93F",X"FB12",X"06F7",X"061D",X"1455",
		X"177B",X"15E1",X"1FA0",X"1EC2",X"1F4A",X"FB67",X"0265",X"FBD9",X"F683",X"EF8B",X"F280",X"F069",X"F611",X"018F",X"082A",X"1513",
		X"01E7",X"FAB6",X"F331",X"F40B",X"E580",X"EA2C",X"DC0A",X"C8B2",X"C653",X"DB0E",X"D8EB",X"DDC0",X"E7F7",X"EA60",X"EC23",X"EB34",
		X"E774",X"D66C",X"DBAF",X"D9AB",X"C407",X"AFD1",X"C0F3",X"C947",X"D4FA",X"D923",X"EF30",X"FA6B",X"F935",X"0CAD",X"11DC",X"0A57",
		X"0C34",X"006F",X"EDBC",X"E768",X"E6B0",X"EB6C",X"DA6C",X"D686",X"E625",X"F353",X"0036",X"08F5",X"130F",X"19D4",X"135C",X"1FA9",
		X"27FF",X"13E9",X"099D",X"0899",X"FD46",X"F096",X"F463",X"01CB",X"072B",X"0993",X"15ED",X"154F",X"1598",X"18BC",X"1800",X"1726",
		X"06E1",X"F996",X"F81B",X"FDE6",X"0C24",X"10D9",X"12C3",X"1115",X"100E",X"1E30",X"270F",X"1ED8",X"1309",X"1DA8",X"1E53",X"1A0A",
		X"129A",X"0B4A",X"0E8A",X"1813",X"24E6",X"2208",X"1CE7",X"170D",X"186F",X"1409",X"1ACB",X"1A07",X"18CA",X"0EA1",X"0890",X"FD84",
		X"F902",X"065D",X"051D",X"0A4B",X"0178",X"0DE6",X"0B0A",X"12B4",X"2032",X"22AC",X"1B3D",X"1A10",X"133C",X"0789",X"02E7",X"0B08",
		X"15B4",X"FD5C",X"F54E",X"F6E0",X"0342",X"0209",X"FDDA",X"05CE",X"F56E",X"F03A",X"ED37",X"F11B",X"ECD8",X"E4A7",X"E5E0",X"DE89",
		X"E4AD",X"F298",X"F6A7",X"F144",X"EC62",X"EFE4",X"F501",X"F0AB",X"EC10",X"EDAB",X"E3E6",X"DF7C",X"E5F2",X"E6A4",X"E93F",X"DF4E",
		X"DC23",X"DBA2",X"E252",X"E5F9",X"EED4",X"ED8F",X"F09B",X"E8A4",X"F295",X"000D",X"F2CE",X"E635",X"F017",X"EAE0",X"F32E",X"ED3A",
		X"EE50",X"EB1D",X"E19A",X"E722",X"EECE",X"F74A",X"F873",X"005F",X"F44A",X"F1CF",X"EF92",X"09E1",X"FBBD",X"F6FC",X"F493",X"FA0C",
		X"F6C0",X"FC4C",X"0469",X"01F0",X"FD2F",X"F919",X"01E4",X"0097",X"0EBA",X"18EB",X"1515",X"07B6",X"0EDF",X"18EE",X"1F31",X"1DDC",
		X"18ED",X"083D",X"04FD",X"0EB7",X"149B",X"123B",X"0C1E",X"028B",X"FC2C",X"00CD",X"0815",X"090E",X"0A9A",X"0CD6",X"091E",X"166C",
		X"1752",X"1E96",X"1DEE",X"22D2",X"2283",X"175C",X"1313",X"10BA",X"0DF5",X"0D2C",X"1191",X"1497",X"1171",X"085A",X"0C54",X"12DC",
		X"1042",X"0890",X"0C84",X"0B51",X"F905",X"F75A",X"FE0D",X"F602",X"F246",X"F5DB",X"FAFC",X"EFC5",X"F7B3",X"0F0B",X"0B1F",X"0B1A",
		X"2867",X"2E68",X"140F",X"0756",X"1358",X"178E",X"FE71",X"FBD6",X"0172",X"F605",X"F28B",X"0550",X"1136",X"1065",X"0F94",X"1216",
		X"11C4",X"0B18",X"120F",X"0C8A",X"FDD6",X"F4F2",X"F344",X"F4E8",X"EFE2",X"ED14",X"F1CE",X"E26A",X"EEFD",X"F8A9",X"F007",X"F734",
		X"F24E",X"E5B3",X"DF44",X"E322",X"EB65",X"EFFB",X"F26A",X"F550",X"ECCD",X"F217",X"002C",X"F7F5",X"F841",X"E1A7",X"D5B4",X"BC55",
		X"B5FC",X"BC29",X"D4B1",X"E365",X"D776",X"DB5C",X"D552",X"F602",X"121F",X"2587",X"1EB6",X"1613",X"13AA",X"0DF3",X"FFDA",X"FB5B",
		X"F1B9",X"D546",X"C214",X"CA46",X"E5A7",X"FCDD",X"0990",X"0A41",X"0DD6",X"1E41",X"3573",X"2EF1",X"193A",X"0B02",X"0A27",X"0424",
		X"F527",X"F71B",X"FEC9",X"FA12",X"FD61",X"0E8D",X"1E01",X"25B6",X"2A91",X"39E2",X"3BBD",X"2EB2",X"1406",X"10B7",X"0502",X"01C4",
		X"04D1",X"09E8",X"0CEB",X"0F15",X"1119",X"207D",X"1749",X"11E9",X"22D9",X"203E",X"126B",X"0CFC",X"11E0",X"09A6",X"F2CF",X"F341",
		X"025F",X"0042",X"0DB9",X"1300",X"1B99",X"0E58",X"1067",X"0FD7",X"18E7",X"0A05",X"0876",X"08B9",X"FC65",X"EE8C",X"F48C",X"01AE",
		X"FF3F",X"0262",X"15B0",X"13A1",X"0085",X"0D76",X"0D4B",X"0F7E",X"FE35",X"FC06",X"EBDA",X"DEC2",X"F22A",X"0B99",X"0EC9",X"FF72",
		X"FFE0",X"F8DC",X"EC4C",X"DD01",X"E390",X"E199",X"D68B",X"D094",X"D1F3",X"ECAC",X"029E",X"11DA",X"1041",X"11E7",X"0B67",X"06E2",
		X"02F4",X"0279",X"FB71",X"E4BD",X"CCBC",X"BAD7",X"B454",X"C49C",X"CC22",X"D0C1",X"D2A7",X"E3F6",X"FF53",X"0A25",X"1148",X"1F2E",
		X"1939",X"0796",X"0C1E",X"0C57",X"FC06",X"DCB6",X"CA83",X"C050",X"BC5B",X"D041",X"FFFC",X"09C5",X"077F",X"12BD",X"1E80",X"1E8A",
		X"102B",X"1510",X"FF2F",X"E0DD",X"E96C",X"F89A",X"F3CC",X"E88E",X"F06F",X"0489",X"FD7B",X"F96D",X"F4CF",X"FAC0",X"0036",X"09DE",
		X"1A1A",X"18E8",X"0D22",X"0880",X"0B5E",X"EF9E",X"F463",X"F311",X"F744",X"F10E",X"FA84",X"0146",X"FE39",X"0546",X"1752",X"1901",
		X"0F4B",X"1C2A",X"16B8",X"0F45",X"0F18",X"1A53",X"1064",X"0082",X"F9FB",X"07D2",X"0EA6",X"1105",X"1746",X"250E",X"2712",X"1E54",
		X"0ED9",X"0333",X"FCDC",X"00E3",X"FEEE",X"0346",X"048B",X"107B",X"1C56",X"14F3",X"0E06",X"0F13",X"2654",X"28D7",X"1F15",X"20B6",
		X"2212",X"1CC2",X"120C",X"1CF1",X"29C7",X"1E60",X"1D6D",X"1665",X"0611",X"EC21",X"ECF3",X"EC6C",X"E6CD",X"E419",X"F4EC",X"050B",
		X"0C28",X"0B54",X"1D43",X"222B",X"19A5",X"19AB",X"0A54",X"037F",X"05E2",X"0BA3",X"FBC7",X"F89A",X"EF20",X"EA82",X"FB45",X"0CD6",
		X"083D",X"0CBC",X"1125",X"20BF",X"1ADA",X"169A",X"16FE",X"126E",X"039B",X"FD03",X"08AA",X"0663",X"06D1",X"FC25",X"0867",X"0450",
		X"0EF9",X"2F52",X"3B44",X"2BD3",X"2028",X"2C3F",X"2F50",X"1E5C",X"1CD4",X"2105",X"096A",X"02A5",X"1D2A",X"1DBC",X"169E",X"2635",
		X"28AA",X"1623",X"0292",X"26F6",X"1D53",X"08B3",X"0AD2",X"0D05",X"0AA6",X"0278",X"15BB",X"05F4",X"0AB6",X"14CC",X"1BD2",X"FDED",
		X"025F",X"11CA",X"0DAD",X"051E",X"E9CE",X"E483",X"D7F1",X"DFC3",X"E5F9",X"EA23",X"DDEF",X"D219",X"D859",X"DCF2",X"E1A0",X"E6D0",
		X"F295",X"E406",X"E5CF",X"FBE9",X"048C",X"0D64",X"064D",X"FC7E",X"F440",X"F5C5",X"0676",X"0511",X"FAF0",X"071A",X"0D42",X"0265",
		X"04CD",X"07DC",X"0E87",X"13F6",X"1AD7",X"1226",X"FBC3",X"FDF6",X"FDC7",X"F130",X"ECA5",X"EC62",X"EE13",X"ECB5",X"F2A2",X"FA1B",
		X"FC10",X"FE65",X"018B",X"FCB3",X"FAD7",X"F66A",X"F544",X"EC8B",X"E20F",X"EEDB",X"F3A3",X"E83C",X"EF11",X"03C4",X"0DD3",X"1178",
		X"14ED",X"189E",X"044A",X"0330",X"FFEA",X"ED75",X"DBAF",X"E201",X"E69B",X"EFE8",X"F0D7",X"F0BE",X"EA43",X"EFAF",X"05AF",X"0AC2",
		X"F990",X"F383",X"E8E7",X"E7FC",X"E3F9",X"E084",X"ED23",X"DF05",X"E449",X"E2A0",X"FBE9",X"FAEC",X"0CA9",X"1A2D",X"2412",X"128A",
		X"1985",X"1B50",X"0B8D",X"0EDA",X"097A",X"059E",X"F401",X"0194",X"05E8",X"02CB",X"137F",X"2597",X"3605",X"2919",X"26B1",X"3583",
		X"2A1C",X"2B12",X"2A8E",X"24CC",X"1075",X"09FE",X"1F7D",X"2A33",X"19F4",X"16BA",X"1891",X"142A",X"0DCF",X"0F7D",X"17C8",X"014C",
		X"E88E",X"FADF",X"FF23",X"EC03",X"F4F2",X"0AB9",X"FFCA",X"EE53",X"098A",X"1F1B",X"0B6D",X"F8D9",X"FCB3",X"F84B",X"DEE9",X"EE36",
		X"FBFF",X"E20C",X"D3E7",X"EE46",X"FA6A",X"F673",X"F850",X"0016",X"F221",X"EC62",X"F64D",X"F984",X"E9B1",X"E8B0",X"DF1E",X"E791",
		X"E471",X"ED79",X"FE4F",X"FD7E",X"FDFF",X"FDB4",X"FF65",X"FC8E",X"FE58",X"F140",X"F314",X"D6D7",X"E270",X"DA23",X"D8E7",X"F393",
		X"FE17",X"FFE0",X"F702",X"0744",X"1BA5",X"1749",X"33F4",X"3BF9",X"2089",X"14DD",X"0957",X"FB1C",X"E6CA",X"DB3E",X"E1E0",X"D7AE",
		X"CF94",X"E820",X"ED6F",X"DE9D",X"E002",X"EB36",X"02A5",X"F890",X"F8D6",X"FB77",X"E351",X"E47A",X"01B1",X"0019",X"0120",X"046F",
		X"FBA7",X"F070",X"EF73",X"1358",X"2267",X"1BF1",X"0C1A",X"1FEB",X"1DF7",X"2125",X"2D6C",X"2962",X"0DA3",X"1122",X"1AFD",X"0A0E",
		X"0299",X"034C",X"0869",X"05A9",X"0837",X"093A",X"05E8",X"F6A3",X"F770",X"F615",X"0CF2",X"0B71",X"0986",X"0B08",X"F8E9",X"E484",
		X"F35D",X"134E",X"0DAD",X"FD8B",X"EC76",X"F684",X"F6E9",X"0F5D",X"1E99",X"239A",X"1BAC",X"216D",X"1FF1",X"0F7A",X"F7C2",X"0579",
		X"02D1",X"FA0E",X"E7AA",X"CC80",X"CD11",X"D9D8",X"E8F3",X"E8BA",X"ECD5",X"DD3D",X"E8A4",X"FAD0",X"0F57",X"065D",X"1267",X"1261",
		X"1487",X"11CE",X"155F",X"0F5B",X"1516",X"1D8C",X"1EEF",X"2BD1",X"1F11",X"20B3",X"1F8F",X"25C0",X"2096",X"277E",X"37F8",X"3935",
		X"2E0A",X"25EC",X"1F47",X"0F94",X"0F6E",X"1103",X"092E",X"F7DC",X"FBDC",X"05BB",X"FAA1",X"FBA7",X"08B6",X"0660",X"FB45",X"0398",
		X"0C1B",X"FDE7",X"EA36",X"E819",X"FA5E",X"F37A",X"E393",X"D603",X"C1E4",X"C6E1",X"D5CB",X"EBEA",X"E277",X"DFE2",X"DFF7",X"F1FB",
		X"EFC5",X"F1DE",X"FD32",X"E945",X"E4DA",X"E39D",X"DFAC",X"CEBD",X"C82A",X"CA0A",X"D05C",X"C86A",X"DAA2",X"E7EC",X"ED72",X"F537",
		X"F3C2",X"F217",X"F534",X"EF20",X"FD28",X"F6F2",X"E53C",X"E9F3",X"F8F0",X"0656",X"0072",X"0350",X"0E4F",X"08FE",X"F67D",X"0B30",
		X"FD79",X"FA96",X"0126",X"1090",X"16FA",X"FFCD",X"0B38",X"1D89",X"213A",X"271B",X"2AD7",X"2751",X"120F",X"1C24",X"312D",X"2868",
		X"1746",X"1355",X"1025",X"F6B3",X"F499",X"F247",X"F014",X"DC4A",X"E82F",X"FC38",X"0018",X"0B70",X"0E84",X"1C63",X"1BA2",X"1D3C",
		X"2E03",X"249E",X"1B0A",X"0EC6",X"03D1",X"0905",X"0D83",X"0AFF",X"08E4",X"FA78",X"EA5F",X"E054",X"DF08",X"F633",X"EEC8",X"DAA5",
		X"C2DB",X"BEAA",X"CCFC",X"E231",X"EDCB",X"EA5E",X"E321",X"EBDA",X"06C8",X"0770",X"1E4A",X"2594",X"14CE",X"00FD",X"F2F1",X"077D",
		X"0F85",X"1251",X"0EE6",X"066D",X"017C",X"0AA6",X"06F7",X"0DC3",X"181A",X"1F63",X"23BC",X"2093",X"29E9",X"230C",X"2A45",X"2B1F",
		X"222B",X"17B1",X"18E4",X"0D22",X"00FD",X"FDAD",X"0369",X"0E7D",X"0AF2",X"07CE",X"0CAD",X"FF7B",X"FD69",X"F6C3",X"F8C6",X"083A",
		X"FC75",X"0700",X"EF43",X"ED1C",X"F524",X"09CC",X"0ABB",X"FD2F",X"F5A9",X"E36B",X"D610",X"CE41",X"EC76",X"EA13",X"DF93",X"D578",
		X"D6C7",X"E183",X"F1D8",X"0688",X"0129",X"EE2C",X"FC38",X"0ECC",X"048F",X"ECB1",X"EB5C",X"EBE4",X"F07C",X"F5A3",X"F9D9",X"F4C2",
		X"ECE7",X"EF23",X"FD22",X"0E4B",X"07B2",X"1AF4",X"0C67",X"051A",X"1055",X"28BD",X"2745",X"128F",X"04C8",X"0359",X"EE5D",X"EF75",
		X"07E2",X"FCFA",X"F4D9",X"EFA8",X"F73B",X"05AE",X"FF39",X"0216",X"0162",X"ED96",X"FF00",X"EE0A",X"F7C9",X"F32A",X"EC88",X"E8BB",
		X"F42E",X"EF6A",X"EA4F",X"EEAB",X"F36A",X"FE5C",X"F305",X"0117",X"EEF1",X"F417",X"F7EF",X"E48E",X"DA1A",X"D840",X"E194",X"EB79",
		X"EEBE",X"FDAA",X"0450",X"07F4",X"158E",X"2141",X"24D9",X"3085",X"2099",X"14AE",X"10D5",X"143C",X"1778",X"08F4",X"0027",X"F3AF",
		X"F951",X"0925",X"1AA7",X"1EDB",X"2B3E",X"30D1",X"30EF",X"3E91",X"2842",X"250F",X"21D9",X"0C1A",X"F18D",X"E85C",X"F701",X"ED2C",
		X"FC46",X"0036",X"0B4E",X"022C",X"12F2",X"24D3",X"1F17",X"1AAE",X"0B1F",X"08D5",X"F9BA",X"F9A0",X"09AF",X"0C51",X"F3D6",X"E6AD",
		X"EDFE",X"F637",X"FD2C",X"FC2F",X"FD6B",X"F952",X"EFEB",X"FFE4",X"0C35",X"0867",X"0614",X"1ADB",X"28C6",X"1C75",X"13DA",X"1930",
		X"00FA",X"02BC",X"0834",X"F583",X"DAF1",X"CA9D",X"DB1D",X"EE5C",X"F34A",X"F2FB",X"03B8",X"0A5A",X"18A8",X"259C",X"33AC",X"24D0",
		X"17D4",X"0394",X"FA93",X"F153",X"ED40",X"EFF1",X"DA7C",X"D582",X"DE14",X"FB25",X"0839",X"1210",X"1BC2",X"14E6",X"113C",X"0F67",
		X"16CB",X"FD29",X"DE90",X"E081",X"CF32",X"C8F2",X"C0A2",X"C49C",X"CAC2",X"D01E",X"DD86",X"E61C",X"EC9E",X"EA01",X"EAB5",X"E48D",
		X"DE28",X"DAB6",X"D975",X"D164",X"C963",X"D057",X"D9FE",X"F3BF",X"FC51",X"01AE",X"0FFC",X"0CBF",X"0E3E",X"1328",X"1F2B",X"12A7",
		X"08B6",X"F1A2",X"E518",X"F41E",X"00FD",X"0AC6",X"FFD0",X"F83B",X"F952",X"0082",X"FA3F",X"07B5",X"08EB",X"0227",X"F270",X"EEE7",
		X"0627",X"0578",X"084D",X"11F6",X"1655",X"1351",X"1CDE",X"2C36",X"30F1",X"18CA",X"13B4",X"1B37",X"0459",X"FF6F",X"1142",X"1078",
		X"FE09",X"FC12",X"1A1D",X"25A1",X"220F",X"2B9B",X"27F9",X"1B27",X"21B8",X"2387",X"0BBA",X"F728",X"F282",X"07AF",X"FD3F",X"F8EC",
		X"0566",X"05B8",X"089A",X"139E",X"1A2D",X"1716",X"1C2A",X"20D5",X"15F3",X"03FB",X"0A24",X"127E",X"0659",X"FF48",X"FFB7",X"FD51",
		X"0C51",X"12DD",X"185E",X"0AAF",X"FAD0",X"F83B",X"FDC3",X"0200",X"FEE3",X"F72C",X"F1C8",X"F0D5",X"F2E5",X"05DB",X"08CF",X"FF85",
		X"F3E5",X"F708",X"F1CF",X"FCD3",X"03F3",X"FBC1",X"F62B",X"F9FC",X"05F2",X"02E7",X"05BF",X"01BE",X"F91F",X"EC59",X"F2F2",X"F8CF",
		X"04F1",X"F5BC",X"F296",X"F461",X"0036",X"0F35",X"12B1",X"170A",X"0D05",X"0AFB",X"082A",X"0586",X"F845",X"FCD0",X"0253",X"F06C",
		X"DC53",X"E001",X"EE43",X"E9A1",X"E3E0",X"FE2C",X"F696",X"EEE5",X"0236",X"0C14",X"0401",X"059F",X"F79A",X"E21C",X"DCD8",X"E08E",
		X"EE26",X"DC44",X"CA3E",X"C75A",X"C912",X"DD73",X"EB0A",X"F2D2",X"E72C",X"E608",X"F6FE",X"063A",X"F4A9",X"F7B3",X"F938",X"E312",
		X"D0CD",X"BBFF",X"C48E",X"C7D2",X"D336",X"D9B2",X"DAF5",X"D2E6",X"DF38",X"FD91",X"0D1E",X"FFED",X"FD91",X"FC6E",X"E952",X"F642",
		X"0AAF",X"06BC",X"001D",X"F65A",X"FE16",X"070B",X"09B6",X"115B",X"27D7",X"2FA5",X"2277",X"19DD",X"211A",X"243E",X"236A",X"2E9E",
		X"2BC1",X"213B",X"12E6",X"2322",X"2FA2",X"3296",X"381C",X"3E8B",X"3854",X"2CE6",X"2BC0",X"2A94",X"2A5B",X"20D9",X"2748",X"1FC5",
		X"1792",X"2393",X"221B",X"27C9",X"2FA7",X"3490",X"3D61",X"3C26",X"3289",X"2F9F",X"2D8F",X"30F4",X"1817",X"F9A7",X"0113",X"09D5",
		X"0EA4",X"F977",X"F42B",X"E70D",X"E315",X"E2EF",X"E27D",X"E56E",X"CEA1",X"D9EE",X"D68B",X"DA7C",X"EAD4",X"FD38",X"0AAC",X"F5E2",
		X"E8A4",X"F48D",X"0323",X"031D",X"01FA",X"E9AE",X"D085",X"C026",X"C7DC",X"E0A0",X"DF07",X"E31F",X"DBE7",X"E615",X"E9A7",X"F6FF",
		X"0488",X"080B",X"0D6E",X"F9E8",X"F108",X"EC6C",X"F951",X"FCA7",X"0592",X"05EB",X"F928",X"EFCB",X"FD3C",X"0006",X"F62B",X"FB32",
		X"F40B",X"EADA",X"E2C3",X"FCAA",X"0686",X"0E35",X"0BEF",X"1917",X"188C",X"14E0",X"20DC",X"24C0",X"10AE",X"F076",X"F273",X"EBF1",
		X"DA96",X"C724",X"CD51",X"CA15",X"D287",X"E03E",X"FC68",X"0931",X"1519",X"15D7",X"0BE9",X"11E7",X"1071",X"00F7",X"EE2A",X"E0AD",
		X"E5BD",X"E23E",X"CDC3",X"D131",X"D4D7",X"E1D8",X"F944",X"0D54",X"0863",X"05A6",X"FE40",X"093D",X"0255",X"047F",X"F192",X"D54C",
		X"C89F",X"DF46",X"F7C5",X"F631",X"0860",X"1609",X"161A",X"113F",X"2DFD",X"31EB",X"1EA8",X"0E87",X"153F",X"0D32",X"FFFF",X"FF1A",
		X"FF4F",X"E765",X"EB2A",X"F76B",X"F166",X"EFE7",X"FBA4",X"FE35",X"EDB2",X"F269",X"15C7",X"2102",X"0CB8",X"0BAD",X"1552",X"236E",
		X"1DF5",X"294F",X"2D1A",X"25BD",X"18E4",X"146F",X"0960",X"F645",X"1258",X"1655",X"1297",X"0598",X"1636",X"1E99",X"1297",X"20BD",
		X"2AC7",X"1FD2",X"094A",X"070E",X"07AB",X"0042",X"FEE4",X"0DD3",X"02ED",X"0B05",X"0A21",X"1A39",X"21E5",X"207A",X"2A3C",X"2B1A",
		X"3369",X"3728",X"193A",X"128E",X"0D44",X"01F7",X"FD7B",X"FD52",X"06BC",X"FDE6",X"FA29",X"0E67",X"10C9",X"2209",X"2D65",X"1C14",
		X"0EAC",X"0424",X"0DA9",X"F7B2",X"E8FA",X"DE30",X"D5F6",X"C23D",X"C06C",X"C580",X"D426",X"D3CE",X"E0A0",X"F0DB",X"F75A",X"FADC",
		X"F3B6",X"ECCD",X"EA92",X"F24A",X"ED3D",X"DF6A",X"D34C",X"DBBB",X"D306",X"CD47",X"D4A8",X"D5C7",X"D129",X"DA9F",X"EA17",X"F566",
		X"E1F4",X"DC60",X"F725",X"EF92",X"E50F",X"E2D0",X"DCC8",X"D820",X"E325",X"FB91",X"0AE8",X"003F",X"0B83",X"1AD4",X"0BDE",X"FED9",
		X"12CA",X"2B6B",X"1672",X"072A",X"0617",X"0B21",X"F711",X"FCC7",X"07AF",X"F2B8",X"E157",X"E6CD",X"F6CC",X"F87E",X"FEEB",X"0C61",
		X"0A51",X"FE06",X"FB1C",X"1888",X"2887",X"0DAA",X"0D6E",X"06D8",X"FC64",X"EF7C",X"F928",X"FFED",X"EBAF",X"CF4B",X"DE66",X"E8E7",
		X"EAA4",X"F7A3",X"FA03",X"F8F6",X"EBCB",X"FAF2",X"1247",X"0E3E",X"0C05",X"10C9",X"0EE3",X"0B2B",X"05CF",X"1733",X"161C",X"0620",
		X"014F",X"19D4",X"1823",X"196F",X"2694",X"3E2C",X"2CE4",X"2AE1",X"3EE1",X"248D",X"1297",X"187F",X"1C66",X"0DC0",X"FAF9",X"0617",
		X"0F24",X"FDC0",X"167E",X"2616",X"2D69",X"19FD",X"2AC0",X"3A94",X"262F",X"1F3E",X"2761",X"256E",X"1636",X"0EB7",X"0C34",X"0534",
		X"F501",X"FD0F",X"FFBB",X"FBF6",X"01DE",X"08FB",X"0A80",X"F89A",X"FB52",X"145B",X"1019",X"04E2",X"F86B",X"DC18",X"DAC8",X"E75B",
		X"E681",X"E5CD",X"D8A9",X"D86F",X"D9A5",X"E471",X"F518",X"FAE0",X"EFE8",X"F073",X"EC00",X"EF85",X"EBCE",X"E1CF",X"E55F",X"D8A8",
		X"E0F1",X"E859",X"ED75",X"E56B",X"EA69",X"E5C3",X"DFAA",X"ECE4",X"F4E5",X"FD84",X"F68A",X"F505",X"F7FB",X"F9DA",X"0028",X"FFCD",
		X"0416",X"FF2C",X"F11B",X"E122",X"E8C9",X"F1FB",X"EF02",X"F84A",X"F490",X"F2DE",X"EB49",X"F3DB",X"0698",X"08B8",X"0854",X"122E",
		X"1238",X"FE6E",X"F55E",X"09D6",X"138E",X"060E",X"0436",X"F7A6",X"EE82",X"EE63",X"FAF5",X"064A",X"F026",X"ED59",X"FE62",X"FD68",
		X"0772",X"0CEF",X"13FA",X"0967",X"FA19",X"0F08",X"1575",X"FD55",X"0963",X"10EC",X"0FED",X"0D31",X"0656",X"16B5",X"0AE2",X"0B6A",
		X"0A50",X"0386",X"03B5",X"0A80",X"0957",X"01F4",X"EDEE",X"F0AF",X"0210",X"F797",X"0156",X"0D01",X"14BA",X"0E1B",X"0D9D",X"140D",
		X"0DBD",X"16FE",X"1D01",X"1CDE",X"0CCF",X"06EE",X"00FA",X"0510",X"FF58",X"F9DA",X"FBE0",X"E8D3",X"E9D4",X"F453",X"0113",X"0230",
		X"FF71",X"09D8",X"04FA",X"FA5E",X"00F9",X"FE48",X"0793",X"067F",X"08FF",X"0D5D",X"08B5",X"0641",X"085D",X"00AD",X"0356",X"0579",
		X"02DA",X"007B",X"017C",X"0A21",X"FFF0",X"0282",X"0FE3",X"0C67",X"019B",X"FCBA",X"FE45",X"FC13",X"F851",X"FA9A",X"F340",X"EC36",
		X"EC01",X"F957",X"EFF7",X"EC07",X"FFB2",X"13A1",X"0DB9",X"0DB3",X"1EF2",X"1509",X"FE71",X"07BC",X"1DF4",X"1352",X"031D",X"017F",
		X"FCB3",X"F0A5",X"F8D0",X"0890",X"00F6",X"F550",X"FFE7",X"08DB",X"057F",X"007B",X"0B97",X"157B",X"09C5",X"FED7",X"F5B2",X"E39D",
		X"D882",X"D9B8",X"D509",X"D8A2",X"DD28",X"E9D4",X"F0F5",X"EFB2",X"F9FC",X"0844",X"07BF",X"FE71",X"016C",X"FD48",X"FE16",X"F3BF",
		X"F476",X"F42E",X"ED40",X"E612",X"E72F",X"E5E6",X"E6EC",X"EBA7",X"F2B5",X"FBE7",X"FEE6",X"055A",X"077F",X"015C",X"F6AC",X"0092",
		X"FFE7",X"013C",X"FD68",X"FC2F",X"F7D0",X"F773",X"0223",X"0847",X"059F",X"0693",X"0E2F",X"0ED2",X"0EAA",X"1265",X"1998",X"17ED",
		X"135E",X"0EC6",X"09EE",X"FBC6",X"F4DF",X"F5A9",X"FA84",X"022D",X"0BD9",X"0DE6",X"0A66",X"0BEC",X"1BB5",X"24FF",X"1D1E",X"1BFD",
		X"178E",X"1158",X"084D",X"0917",X"0AC9",X"0453",X"FE42",X"F857",X"EF14",X"F096",X"000C",X"0559",X"095F",X"0EA0",X"0F7A",X"138F",
		X"0688",X"0352",X"0401",X"F9C0",X"F941",X"F5E2",X"F6C6",X"F5A3",X"EFE2",X"F247",X"FAEC",X"FF09",X"07BB",X"0478",X"027C",X"01CE",
		X"0546",X"0A8C",X"07AF",X"0062",X"020A",X"FDA7",X"F4E8",X"EF60",X"E49E",X"E3DF",X"E0C8",X"E48D",X"EA13",X"EAE7",X"EEE4",X"F638",
		X"F8E2",X"FF6E",X"0036",X"0BB3",X"102F",X"0235",X"FE72",X"FDE7",X"020A",X"0006",X"FD4B",X"F8F0",X"F317",X"F1F5",X"F4DB",X"FF1C",
		X"FE72",X"048F",X"0245",X"0195",X"070B",X"0D17",X"10C7",X"08BF",X"075A",X"0901",X"0446",X"FA3B",X"F893",X"0029",X"0094",X"FD35",
		X"011D",X"0AA9",X"14EA",X"1556",X"181E",X"18FE",X"169E",X"1400",X"1B31",X"1976",X"1632",X"0A2D",X"004F",X"FA25",X"F997",X"040A",
		X"0550",X"02B8",X"FBA1",X"FE52",X"0621",X"07C1",X"0C14",X"12AA",X"1155",X"0BAC",X"0659",X"08CF",X"0C47",X"0924",X"0376",X"FDCA",
		X"F3F8",X"EC5C",X"EB9E",X"F49A",X"F7F5",X"F51F",X"F75D",X"FB88",X"F9F2",X"F7E2",X"F9A0",X"FA45",X"F694",X"EFB4",X"EB85",X"EA7C",
		X"ED5F",X"F2C2",X"F1BB",X"EF20",X"F1EA",X"F1EB",X"F1F2",X"F247",X"F19E",X"F514",X"F4EB",X"F4FF",X"F6D2",X"F77B",X"F590",X"F5C3",
		X"F39F",X"F0BB",X"F020",X"EE63",X"ED53",X"EF31",X"EF4D",X"EC8F",X"F377",X"F72E",X"FC3E",X"02AD",X"0BCF",X"0D57",X"04C8",X"FF0D",
		X"FF9D",X"FC23",X"FA64",X"F9B3",X"F3E5",X"F108",X"F689",X"FF02",X"FEE6",X"032F",X"0876",X"08A8",X"0413",X"0214",X"02D7",X"03F0",
		X"0540",X"0821",X"0472",X"FDCD",X"FB7B",X"F574",X"F296",X"FC09",X"FFA7",X"FFCA",X"0447",X"09D2",X"1057",X"147E",X"169B",X"147E",
		X"14A7",X"11EC",X"0E51",X"0CBD",X"0CCD",X"0B83",X"0D0C",X"0F0F",X"0FAC",X"0F68",X"12F9",X"12A7",X"0F84",X"13D9",X"16A5",X"15D7",
		X"12AA",X"105B",X"0FD3",X"08EE",X"0692",X"0AE2",X"0AC9",X"0BE6",X"0DD9",X"0F5F",X"0DA3",X"0CEE",X"1102",X"0FC3",X"0BEF",X"0E0F",
		X"0E87",X"0D90",X"0D3C",X"0CCF",X"0917",X"039F",X"FB0C",X"F4A0",X"F095",X"EF5D",X"F007",X"F115",X"F0CB",X"F1DE",X"F60B",X"F790",
		X"F60B",X"F732",X"FB3F",X"FA13",X"F787",X"FA13",X"FE4C",X"FFAA",X"FC12",X"F74D",X"F50F",X"F0D4",X"EC88",X"ED92",X"F0CB",X"F2DE",
		X"F667",X"FA80",X"FEA7",X"FEAE",X"0116",X"FDB7",X"F583",X"F201",X"F441",X"F5A6",X"F5AF",X"F741",X"F8CA",X"FBE0",X"F984",X"F99C",
		X"FBE0",X"FE13",X"0140",X"030F",X"042A",X"0146",X"FD48",X"FC32",X"FE9E",X"0042",X"FD6F",X"FABA",X"FA3F",X"FB09",X"FC00",X"FFAE",
		X"FFBE",X"FC12",X"FADF",X"FCD4",X"FFCD",X"01E7",X"040A",X"0917",X"0885",X"035C",X"0449",X"02ED",X"00D5",X"FE72",X"FBE3",X"F9A0",
		X"F984",X"F8A4",X"F931",X"F931",X"FA06",X"FC06",X"FA5B",X"FBF6",X"FF4C",X"0026",X"FEA1",X"FDDB",X"FD36",X"FE9E",X"FF68",X"FE45",
		X"FB5E",X"F891",X"F663",X"F4BF",X"F55D",X"F9DA",X"FEA4",X"0075",X"0353",X"0524",X"086C",X"08B6",X"080E",X"06A6",X"03A8",X"FF12",
		X"FED3",X"0185",X"035C",X"012A",X"0043",X"020D",X"0345",X"0837",X"087A",X"0847",X"076F",X"06A2",X"07A8",X"0B57",X"092A",X"0808",
		X"03D8",X"028F",X"03AB",X"0200",X"0069",X"FC84",X"FB7E",X"FD0F",X"00A4",X"05F7",X"0947",X"0A7A",X"0B5B",X"0DBD",X"0FE0",X"0D3B",
		X"0BAF",X"0987",X"04B6",X"FEFA",X"FCD9",X"FAC0",X"F7DC",X"F9EC",X"FCC7",X"FC88",X"FCE0",X"FF3C",X"06F5",X"08FF",X"0AA0",X"0F2E",
		X"0F0F",X"0C71",X"0ACC",X"09BC",X"07EF",X"051A",X"00A8",X"FFD1",X"FFDA",X"023D",X"0504",X"05FB",X"074D",X"096F",X"0C96",X"0C18",
		X"0D7E",X"0F67",X"0AF8",X"081B",X"02CB",X"01CB",X"0142",X"FD7B",X"F94F",X"F5C3",X"F705",X"F912",X"FB5E",X"FB96",X"FE6E",X"FF36",
		X"FEBD",X"FB15",X"F9D0",X"FA3E",X"F7FF",X"F5D9",X"F2E8",X"EE6F",X"ED60",X"EBD1",X"EC79",X"EDAE",X"EB89",X"ED52",X"EE5C",X"F180",
		X"F4D9",X"F47D",X"F754",X"F8B3",X"F50B",X"F393",X"F2F5",X"F353",X"F28C",X"EF5A",X"EE56",X"ECC5",X"ECA8",X"F1EC",X"F35A",X"F440",
		X"F59A",X"FA9D",X"FB91",X"FA2B",X"FC78",X"FECA",X"FE71",X"FD0C",X"FD39",X"FD81",X"FCA7",X"FAF2",X"FE29",X"0026",X"FF5B",X"FFA1",
		X"025C",X"03BF",X"0365",X"06BC",X"093D",X"0C35",X"0E6B",X"0BE6",X"0B48",X"0D28",X"0F97",X"0CA6",X"060B",X"049B",X"03E7",X"0330",
		X"05EE",X"0801",X"098A",X"0A20",X"0D37",X"0DEE",X"0D3F",X"109D",X"1422",X"155C",X"13FA",X"0DD9",X"08F1",X"0411",X"FF26",X"FD61",
		X"FA38",X"F8C2",X"F915",X"F968",X"FAEC",X"024A",X"07E5",X"0A92",X"0AE9",X"09D2",X"0B9F",X"0BC3",X"0A01",X"069E",X"00EA"
	);
begin
	process(clk)
	begin
		if rising_edge(clk) then
			if addr=x"ffff" then
				data <= (others => '0');
			else
				data <= rom_data(to_integer(unsigned(addr)));
			end if;
		end if;
	end process;
end architecture;
